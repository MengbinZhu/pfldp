netcdf ropp_test_2v {
dimensions:
	dim_unlim = UNLIMITED ; // (1 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1a = 100 ;
	dim_lev1b = 100 ;
	dim_lev2a = 100 ;
	dim_lev2b = 100 ;
	dim_lev2d = 100 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 360. ;
	char bg_source(dim_unlim, dim_char20) ;
		bg_source:long_name = "Background data source" ;
	int bg_year(dim_unlim) ;
		bg_year:long_name = "VT year" ;
		bg_year:units = "years" ;
		bg_year:valid_range = 1995, 2099 ;
	int bg_month(dim_unlim) ;
		bg_month:long_name = "VT month" ;
		bg_month:units = "months" ;
		bg_month:valid_range = 1, 12 ;
	int bg_day(dim_unlim) ;
		bg_day:long_name = "VT day" ;
		bg_day:units = "days" ;
		bg_day:valid_range = 1, 31 ;
	int bg_hour(dim_unlim) ;
		bg_hour:long_name = "VT hour" ;
		bg_hour:units = "hours" ;
		bg_hour:valid_range = 0, 23 ;
	int bg_minute(dim_unlim) ;
		bg_minute:long_name = "VT minute" ;
		bg_minute:units = "minutes" ;
		bg_minute:valid_range = 0, 59 ;
	float bg_fcperiod(dim_unlim) ;
		bg_fcperiod:long_name = "Forecast period" ;
		bg_fcperiod:units = "hours" ;
		bg_fcperiod:valid_range = 0., 24. ;
	double dtime(dim_unlim, dim_lev1a) ;
		dtime:long_name = "Time since start of occultation" ;
		dtime:units = "seconds" ;
		dtime:valid_range = -1., 240. ;
	float snr_L1ca(dim_unlim, dim_lev1a) ;
		snr_L1ca:long_name = "Signal-to-noise ratio (L1, C/A code)" ;
		snr_L1ca:units = "volt / volt" ;
		snr_L1ca:valid_range = 0., 50000. ;
	float snr_L1p(dim_unlim, dim_lev1a) ;
		snr_L1p:long_name = "Signal-to-noise ratio (L1, P code)" ;
		snr_L1p:units = "volt / volt" ;
		snr_L1p:valid_range = 0., 50000. ;
	float snr_L2p(dim_unlim, dim_lev1a) ;
		snr_L2p:long_name = "Signal-to-noise ratio (L2, P code)" ;
		snr_L2p:units = "volt / volt" ;
		snr_L2p:valid_range = 0., 50000. ;
	double phase_L1(dim_unlim, dim_lev1a) ;
		phase_L1:long_name = "Excess phase (L1)" ;
		phase_L1:units = "metres" ;
		phase_L1:valid_range = -1.e+06, 1.e+06 ;
	double phase_L2(dim_unlim, dim_lev1a) ;
		phase_L2:long_name = "Excess phase (L2)" ;
		phase_L2:units = "metres" ;
		phase_L2:valid_range = -1.e+06, 1.e+06 ;
	double r_gns(dim_unlim, xyz, dim_lev1a) ;
		r_gns:long_name = "GNSS transmitter position" ;
		r_gns:units = "metres" ;
		r_gns:valid_range = -4.3e+07, 4.3e+07 ;
		r_gns:reference_frame = "ECF" ;
	double v_gns(dim_unlim, xyz, dim_lev1a) ;
		v_gns:long_name = "GNSS transmitter velocity" ;
		v_gns:units = "metres / seconds" ;
		v_gns:valid_range = -10000., 10000. ;
		v_gns:reference_frame = "ECI" ;
	double r_leo(dim_unlim, xyz, dim_lev1a) ;
		r_leo:long_name = "LEO transmitter position" ;
		r_leo:units = "metres" ;
		r_leo:valid_range = -1.e+07, 1.e+07 ;
		r_leo:reference_frame = "ECF" ;
	double v_leo(dim_unlim, xyz, dim_lev1a) ;
		v_leo:long_name = "LEO transmitter velocity" ;
		v_leo:units = "metres / seconds" ;
		v_leo:valid_range = -10000., 10000. ;
		v_leo:reference_frame = "ECI" ;
	float phase_qual(dim_unlim, dim_lev1a) ;
		phase_qual:long_name = "Quality value for phase (and SNR)" ;
		phase_qual:units = "percent" ;
		phase_qual:valid_range = 0., 100. ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 360. ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float alt_refrac(dim_unlim, dim_lev2a) ;
		alt_refrac:long_name = "Geometric height above geoid for refractivity" ;
		alt_refrac:units = "metres" ;
		alt_refrac:valid_range = -1000., 1.e+05 ;
	float geop_refrac(dim_unlim, dim_lev2a) ;
		geop_refrac:long_name = "Geopotential height above geoid for refractivity" ;
		geop_refrac:units = "geopotential metres" ;
		geop_refrac:valid_range = -1000., 1.e+05 ;
	double refrac(dim_unlim, dim_lev2a) ;
		refrac:long_name = "Refractivity" ;
		refrac:units = "N-units" ;
		refrac:valid_range = 0., 500. ;
	double refrac_sigma(dim_unlim, dim_lev2a) ;
		refrac_sigma:long_name = "Estimated error (1-sigma) for refractivity" ;
		refrac_sigma:units = "N-units" ;
		refrac_sigma:valid_range = 0., 50. ;
	float refrac_qual(dim_unlim, dim_lev2a) ;
		refrac_qual:long_name = "Quality value for refractivity" ;
		refrac_qual:units = "percent" ;
		refrac_qual:valid_range = 0., 100. ;
	double dry_temp(dim_unlim, dim_lev2a) ;
		dry_temp:long_name = "Dry temperature" ;
		dry_temp:units = "kelvin" ;
		dry_temp:valid_range = 150., 350. ;
	double dry_temp_sigma(dim_unlim, dim_lev2a) ;
		dry_temp_sigma:long_name = "Estimated error (1-sigma) for dry temperature" ;
		dry_temp_sigma:units = "kelvin" ;
		dry_temp_sigma:valid_range = 0., 50. ;
	float dry_temp_qual(dim_unlim, dim_lev2a) ;
		dry_temp_qual:long_name = "Quality value for dry temperature" ;
		dry_temp_qual:units = "percent" ;
		dry_temp_qual:valid_range = 0., 100. ;
	float geop(dim_unlim, dim_lev2b) ;
		geop:long_name = "Geopotential height above geoid for P,T,H" ;
		geop:units = "geopotential metres" ;
		geop:valid_range = -1000., 1.e+05 ;
	float geop_sigma(dim_unlim, dim_lev2b) ;
		geop_sigma:long_name = "Estimated error (1-sigma) for geopotential height" ;
		geop_sigma:units = "geopotential metres" ;
		geop_sigma:valid_range = 0., 500. ;
	double press(dim_unlim, dim_lev2b) ;
		press:long_name = "Pressure" ;
		press:units = "hPa" ;
		press:valid_range = 0.0001, 1100. ;
	float press_sigma(dim_unlim, dim_lev2b) ;
		press_sigma:long_name = "Estimated error (1-sigma) for pressure" ;
		press_sigma:units = "hPa" ;
		press_sigma:valid_range = 0., 5. ;
	double temp(dim_unlim, dim_lev2b) ;
		temp:long_name = "Temperature" ;
		temp:units = "kelvin" ;
		temp:valid_range = 150., 350. ;
	float temp_sigma(dim_unlim, dim_lev2b) ;
		temp_sigma:long_name = "Estimated error (1-sigma) for temperature" ;
		temp_sigma:units = "kelvin" ;
		temp_sigma:valid_range = 0., 5. ;
	double shum(dim_unlim, dim_lev2b) ;
		shum:long_name = "Specific humidity" ;
		shum:units = "gram / kilogram" ;
		shum:valid_range = 0., 50. ;
	float shum_sigma(dim_unlim, dim_lev2b) ;
		shum_sigma:long_name = "Estimated  error (1-sigma) in specific humidity" ;
		shum_sigma:units = "gram / kilogram" ;
		shum_sigma:valid_range = 0., 5. ;
	float meteo_qual(dim_unlim, dim_lev2b) ;
		meteo_qual:long_name = "Quality value for meteorological data" ;
		meteo_qual:units = "percent" ;
		meteo_qual:valid_range = 0., 100. ;
	float geop_sfc(dim_unlim) ;
		geop_sfc:long_name = "Surface geopotential height" ;
		geop_sfc:units = "geopotential metres" ;
		geop_sfc:valid_range = -1000., 10000. ;
	float press_sfc(dim_unlim) ;
		press_sfc:long_name = "Surface pressure" ;
		press_sfc:units = "hPa" ;
		press_sfc:valid_range = 250., 1100. ;
	float press_sfc_sigma(dim_unlim) ;
		press_sfc_sigma:long_name = "Estimated error (1-sigma) for surface pressure" ;
		press_sfc_sigma:units = "hPa" ;
		press_sfc_sigma:valid_range = 0., 5. ;
	float press_sfc_qual(dim_unlim) ;
		press_sfc_qual:long_name = "Surface pressure quality value" ;
		press_sfc_qual:units = "percent" ;
		press_sfc_qual:valid_range = 0., 100. ;
	double tph_bangle(dim_unlim) ;
		tph_bangle:long_name = "Bending angle-based TPH" ;
		tph_bangle:units = "metres" ;
		tph_bangle:valid_range = 6.2e+06, 6.6e+06 ;
	double tpa_bangle(dim_unlim) ;
		tpa_bangle:long_name = "Bending angle-based TPA" ;
		tpa_bangle:units = "radians" ;
		tpa_bangle:valid_range = -0.001, 0.1 ;
	int tph_bangle_flag(dim_unlim) ;
		tph_bangle_flag:long_name = "Bending angle-based TPH QC flag" ;
		tph_bangle_flag:units = "1" ;
		tph_bangle_flag:valid_range = 0, 255 ;
	float tph_refrac(dim_unlim) ;
		tph_refrac:long_name = "Refractivity-based TPH" ;
		tph_refrac:units = "metres" ;
		tph_refrac:valid_range = -1000., 1.e+05 ;
	double tpn_refrac(dim_unlim) ;
		tpn_refrac:long_name = "Refractivity-based TPN" ;
		tpn_refrac:units = "N-units" ;
		tpn_refrac:valid_range = 0., 500. ;
	int tph_refrac_flag(dim_unlim) ;
		tph_refrac_flag:long_name = "Refractivity-based TPH QC flag" ;
		tph_refrac_flag:units = "1" ;
		tph_refrac_flag:valid_range = 0, 255 ;
	float tph_tdry_lrt(dim_unlim) ;
		tph_tdry_lrt:long_name = "Dry temperature-based TPH (lapse rate)" ;
		tph_tdry_lrt:units = "metres" ;
		tph_tdry_lrt:valid_range = -1000., 1.e+05 ;
	float tpt_tdry_lrt(dim_unlim) ;
		tpt_tdry_lrt:long_name = "Dry temperature-based TPT (lapse rate)" ;
		tpt_tdry_lrt:units = "kelvin" ;
		tpt_tdry_lrt:valid_range = 150., 350. ;
	int tph_tdry_lrt_flag(dim_unlim) ;
		tph_tdry_lrt_flag:long_name = "Dry temperature-based TPH QC flag (lapse rate)" ;
		tph_tdry_lrt_flag:units = "1" ;
		tph_tdry_lrt_flag:valid_range = 0, 255 ;
	float tph_tdry_cpt(dim_unlim) ;
		tph_tdry_cpt:long_name = "Dry temperature-based TPH (cold point)" ;
		tph_tdry_cpt:units = "metres" ;
		tph_tdry_cpt:valid_range = -1000., 1.e+05 ;
	float tpt_tdry_cpt(dim_unlim) ;
		tpt_tdry_cpt:long_name = "Dry temperature-based TPT (cold point)" ;
		tpt_tdry_cpt:units = "kelvin" ;
		tpt_tdry_cpt:valid_range = 150., 350. ;
	int tph_tdry_cpt_flag(dim_unlim) ;
		tph_tdry_cpt_flag:long_name = "Dry temperature-based TPH QC flag (cold point)" ;
		tph_tdry_cpt_flag:units = "1" ;
		tph_tdry_cpt_flag:valid_range = 0, 255 ;
	float prh_tdry_cpt(dim_unlim) ;
		prh_tdry_cpt:long_name = "Dry temperature-based PRH (cold point)" ;
		prh_tdry_cpt:units = "metres" ;
	float prt_tdry_cpt(dim_unlim) ;
		prt_tdry_cpt:long_name = "Dry temperature-based PRT (cold point)" ;
		prt_tdry_cpt:units = "kelvin" ;
	int prh_tdry_cpt_flag(dim_unlim) ;
		prh_tdry_cpt_flag:long_name = "Dry temperature-based PRH QC flag (cold point)" ;
		prh_tdry_cpt_flag:units = "1" ;
	float tph_temp_lrt(dim_unlim) ;
		tph_temp_lrt:long_name = "Temperature-based TPH (lapse rate)" ;
		tph_temp_lrt:units = "geopotential metres" ;
		tph_temp_lrt:valid_range = -1000., 1.e+05 ;
	float tpt_temp_lrt(dim_unlim) ;
		tpt_temp_lrt:long_name = "Temperature-based TPT (lapse rate)" ;
		tpt_temp_lrt:units = "kelvin" ;
		tpt_temp_lrt:valid_range = 150., 350. ;
	int tph_temp_lrt_flag(dim_unlim) ;
		tph_temp_lrt_flag:long_name = "Temperature-based TPH QC flag (lapse rate)" ;
		tph_temp_lrt_flag:units = "1" ;
		tph_temp_lrt_flag:valid_range = 0, 255 ;
	float tph_temp_cpt(dim_unlim) ;
		tph_temp_cpt:long_name = "Temperature-based TPH (cold point)" ;
		tph_temp_cpt:units = "geopotential metres" ;
		tph_temp_cpt:valid_range = -1000., 1.e+05 ;
	float tpt_temp_cpt(dim_unlim) ;
		tpt_temp_cpt:long_name = "Temperature-based TPT (cold point)" ;
		tpt_temp_cpt:units = "kelvin" ;
		tpt_temp_cpt:valid_range = 150., 350. ;
	int tph_temp_cpt_flag(dim_unlim) ;
		tph_temp_cpt_flag:long_name = "Temperature-based TPH QC flag (cold point)" ;
		tph_temp_cpt_flag:units = "1" ;
		tph_temp_cpt_flag:valid_range = 0, 255 ;
	float prh_temp_cpt(dim_unlim) ;
		prh_temp_cpt:long_name = "Temperature-based PRH (cold point)" ;
		prh_temp_cpt:units = "metres" ;
	float prt_temp_cpt(dim_unlim) ;
		prt_temp_cpt:long_name = "Temperature-based PRT (cold point)" ;
		prt_temp_cpt:units = "kelvin" ;
	int prh_temp_cpt_flag(dim_unlim) ;
		prh_temp_cpt_flag:long_name = "Temperature-based PRH QC flag (cold point)" ;
		prh_temp_cpt_flag:units = "1" ;
	char level_type(dim_unlim, dim_char64) ;
		level_type:long_name = "Vertical level type" ;
	float level_coeff_a(dim_unlim, dim_lev2d) ;
		level_coeff_a:long_name = "Hybrid / Eta level coefficient (a or eta)" ;
		level_coeff_a:units = "hPa" ;
		level_coeff_a:valid_range = 0., 2000. ;
	float level_coeff_b(dim_unlim, dim_lev2d) ;
		level_coeff_b:long_name = "Hybrid / Eta level coefficient (b or tau)" ;
		level_coeff_b:units = "1" ;
		level_coeff_b:valid_range = 0., 2. ;

// global attributes:
		:title = "Atmospheric background data for ROPP Radio Occultation data" ;
		:institution = "METO" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "UCAR" ;
		:processing_date = "2014-11-28 14:34:44.196" ;
		:pod_method = "POD_3" ;
		:phase_method = "PHASE_5" ;
		:bangle_method = "BANGLE_2" ;
		:refrac_method = "REFRAC_3" ;
		:meteo_method = "T-DRY" ;
		:thin_method = "SGLIN" ;
		:software_version = "V96.033" ;
		:_FillValue = -9.9999e+07 ;
data:

 occ_id =
  "BG_20141112212842_CO03_R012_UCAR" ;

 gns_id =
  "R012" ;

 leo_id =
  "CO03" ;

 stn_id =
  "PADO" ;

 start_time = 4.6914e+08 ;

 year = 2014 ;

 month = 11 ;

 day = 12 ;

 hour = 21 ;

 minute = 28 ;

 second = 42 ;

 msec = 856 ;

 pcd = 29873 ;

 overall_qual = 4.9989 ;

 time = 4.6914e+08 ;

 time_offset = 106.93 ;

 lat = 53.721 ;

 lon = 172.34 ;

 undulation = 86.256 ;

 roc = 6.2294e+06 ;

 r_coc =
  -14445, -20745, -6612 ;

 azimuth = 138.31 ;

 bg_source =
  "METO" ;

 bg_year = 2014 ;

 bg_month = 11 ;

 bg_day = 12 ;

 bg_hour = 1 ;

 bg_minute = 0 ;

 bg_fcperiod = 13 ;

 dtime =
  25.994, 231.05, 27.347, 100.52, 146.9, 83.477, 84.257, 185.2, 58.956, 
    115.33, 69.08, 125.66, 40.358, 134.93, 220.9, 107.01, 210.56, 48.862, 
    164.84, 137.54, 37.297, 151.1, 52.806, 225.28, 78.287, 12.236, 101.28, 
    191.15, 49.812, 23.767, 109.67, 178.07, 190.45, 202.87, 20.931, 22.979, 
    93.723, 36.536, 24.411, 158.08, 62.264, 2.339, 185.74, 156.08, 140.78, 
    183.18, 50.003, 100.67, 71.337, 133.92, 188.74, 70.336, 116.42, 115.66, 
    118.37, 137.21, 191.06, 228.87, 130.77, 25.126, 122.44, 75.254, 96.834, 
    5.1105, 120.05, 158.36, 46.519, 45.164, 233.19, 83.619, 130.69, 6.9515, 
    11.311, 163.2, 70.661, 122.72, 186.78, 105.68, 24.489, 129.86, 207.73, 
    83.164, 145.16, 33.19, 162.27, 105.74, 198.04, 185.07, 184.2, 208.99, 
    116.74, 24.675, 41.58, 158.34, 42.445, 112.33, 189.04, 38.371, 215.25, 
    112.28 ;

 snr_L1ca =
  17453, 23927, 23040, 27659, 44317, 16694, 9883.3, 26646, 15234, 23697, 
    28573, 43455, 4783.8, 7794.5, 37587, 32619, 33556, 8323.2, 33681, 46306, 
    25845, 18694, 39531, 1548.4, 7624.5, 40689, 43397, 15755, 46891, 18331, 
    47923, 4825.6, 17570, 32949, 47044, 43812, 42745, 36374, 7869.2, 46264, 
    7093.3, 739.34, 20805, 4096.3, 39372, 28023, 34913, 27414, 11289, 29298, 
    6016.2, 18532, 40408, 8541.4, 933.79, 46487, 16948, 7450.8, 36352, 28996, 
    36133, 24094, 38508, 29089, 7983, 20466, 20335, 26935, 14248, 11293, 
    33563, 8615.6, 47088, 4696.8, 22036, 14506, 46611, 40595, 32307, 30273, 
    29243, 6785.9, 22834, 10777, 38353, 37523, 46027, 14826, 24927, 20990, 
    30072, 38053, 46550, 43190, 32658, 14472, 4645.3, 2559, 26149, 29568 ;

 snr_L1p =
  45247, 40790, 27757, 21433, 4681.3, 42257, 47423, 41169, 11626, 6971.9, 
    46149, 18112, 28386, 35257, 19552, 6583.1, 43988, 29979, 12737, 3635.2, 
    43872, 24141, 46719, 41126, 47373, 42936, 8304.4, 39261, 7019.1, 2526.7, 
    41448, 31016, 19449, 3296.1, 41842, 26010, 20008, 35981, 17352, 438.97, 
    33643, 8270.3, 12992, 18634, 10089, 3416.4, 1357.2, 1921.8, 48396, 14647, 
    9728.9, 30555, 42935, 46124, 27701, 20806, 38389, 38870, 35294, 40278, 
    34779, 3446.2, 7026.4, 43939, 34153, 30929, 22352, 5992.3, 13880, 10313, 
    7798.8, 25234, 36997, 19650, 1849.3, 384.3, 6700, 25644, 16488, 8791.1, 
    13963, 45802, 29105, 48207, 6374.9, 23513, 7723.8, 37140, 7190.7, 27379, 
    8933.6, 9637.2, 32135, 19067, 28806, 15180, 14649, 17961, 34947, 40291 ;

 snr_L2p =
  5296.3, 42214, 9478.8, 27672, 8414.2, 48692, 14221, 39146, 47040, 24685, 
    11706, 38217, 24298, 3005.3, 4514.6, 31422, 12760, 8780.8, 3850.4, 40198, 
    31672, 28818, 16276, 6193.3, 47427, 21954, 34521, 11583, 31553, 35873, 
    19.821, 27161, 10537, 7424.4, 22069, 45097, 41452, 1963.4, 15964, 24531, 
    17803, 21146, 7613, 312.62, 1599.6, 20776, 45077, 3501.2, 24005, 36819, 
    17889, 22604, 31118, 5499.2, 46564, 39245, 22392, 18692, 11496, 28931, 
    24224, 17865, 39554, 33638, 32181, 16798, 36007, 45478, 11760, 5484, 
    15396, 19356, 23331, 45083, 11127, 163.04, 39672, 2129.2, 10465, 10694, 
    22388, 41546, 14324, 37554, 48149, 11888, 43694, 34865, 29076, 32239, 
    45037, 43037, 38359, 45689, 4602.6, 19141, 35336, 5736.6, 45630, 25730 ;

 phase_L1 =
  -67950, 8.4951e+05, -4.9513e+05, -2.7784e+05, 8.3045e+05, -3.0814e+05, 
    9.1731e+05, -3.2244e+05, -6.7074e+05, -9.9764e+05, -2.1388e+05, 
    7.6017e+05, -5.8812e+05, -6.6123e+05, 5.1035e+05, 5.467e+05, 5.3156e+05, 
    -62087, 8.6635e+05, 4.1777e+05, -6.195e+05, -59970, -2.3182e+05, -48178, 
    -9.1291e+05, -4.2124e+05, -3.4754e+05, -8.2408e+05, 3.7562e+05, 
    2.082e+05, -4.5629e+05, -4.7946e+05, -3.2512e+05, -1.3778e+05, 
    -3.1515e+05, -1.3747e+05, -8.6777e+05, -8.351e+05, 1.5352e+05, 
    5.0794e+05, -6.3708e+05, -4.5335e+05, 3.3288e+05, -9.2654e+05, 
    7.1499e+05, -20832, 2.6042e+05, 5.115e+05, -1.5636e+05, 5.7181e+05, 
    -27158, 3.3791e+05, -2.9835e+05, 1.9711e+05, -6.7447e+05, -9.0376e+05, 
    -5.2107e+05, -7.6498e+05, -4.0841e+05, -2.7312e+05, -2.3688e+05, 
    -3.6293e+05, -9.5653e+05, -22794, 7.8277e+05, 3.6505e+05, 6.9557e+05, 
    8.2136e+05, 1.8612e+05, 4.2969e+05, -2.0007e+05, -6.1185e+05, 7.8547e+05, 
    -2.4383e+05, -6.2721e+05, -2.6964e+05, 3.7564e+05, 8.9964e+05, 
    -3.389e+05, 2.8718e+05, 2.3582e+05, 3.1754e+05, -8.4412e+05, 95984, 
    4.121e+05, -4.7156e+05, 3.5046e+05, 9.4396e+05, 5.6344e+05, 3.9698e+05, 
    7.0577e+05, -4.2005e+05, -9.0529e+05, 7.2022e+05, -8.2731e+05, 
    -7.3633e+05, -8.125e+05, 4.5801e+05, 6.3424e+05, -3.1037e+05 ;

 phase_L2 =
  2.7025e+05, 37968, 4.7964e+05, -5.5553e+05, -5.147e+05, 9.4552e+05, 
    -2.9027e+05, 7.1826e+05, 5.7713e+05, -6.2843e+05, -1.6592e+05, 
    7.8568e+05, 5.5753e+05, -74689, 2.0386e+05, 43625, 3.7747e+05, 
    -3.8762e+05, -7.0272e+05, -7.8382e+05, 3.5942e+05, -9.9441e+05, 
    3.7561e+05, -3.4173e+05, 3.2291e+05, 8.6746e+05, 7.9575e+05, -1.8765e+05, 
    6.5629e+05, 2.4596e+05, 1.1155e+05, -2.7375e+05, -9.0387e+05, 1.2534e+05, 
    9.08e+05, 4.4609e+05, 7.1919e+05, 8.4637e+05, -8.1548e+05, -7.228e+05, 
    5.843e+05, -9.2283e+05, -4.6599e+05, -3.6079e+05, 4.0819e+05, 
    -5.5211e+05, -8.6476e+05, -3.9742e+05, 95790, 5.5338e+05, -5.9932e+05, 
    -4.5134e+05, 3.1868e+05, -49623, 8.1086e+05, 3.8943e+05, 1.6743e+05, 
    59345, -6.7905e+05, -7.3483e+05, 9.1667e+05, 8.9094e+05, 3.0545e+05, 
    -3.6622e+05, 6.3205e+05, -5.1902e+05, 7.8675e+05, 2.2846e+05, 
    -2.9008e+05, -2.2676e+05, 7.862e+05, -4.0385e+05, 3.8993e+05, 
    -1.3552e+05, -3.3251e+05, -3.1063e+05, -7.6807e+05, 4.8076e+05, -69860, 
    -5.2236e+05, 4.44e+05, 1.1879e+05, -59804, 8.3481e+05, 1.7136e+05, 
    -9.8051e+05, 3.9215e+05, 6.5882e+05, -4.776e+05, -2.7879e+05, 8.3098e+05, 
    -7.4217e+05, 7.8218e+05, -2.4605e+05, -6.2289e+05, 7.2417e+05, 1.44e+05, 
    7.2307e+05, -1.8435e+05, -9.2943e+05 ;

 r_gns =
  -2.2607e+06, -2.8784e+07, -8.112e+06, -2.7766e+06, 2.3273e+07, 1.044e+07, 
    8.4441e+05, 9.2184e+06, 1.1871e+07, 4.1491e+06, 1.206e+06, 6.2581e+06, 
    -1.44e+06, -9.7035e+06, -2.4922e+06, -1.6341e+06, -5.8065e+06, 
    3.1172e+06, -2.2297e+07, 3.0751e+07, -1.4378e+07, -7.958e+06, 7.0798e+06, 
    -2.3235e+06, 1.9976e+06, -1.3896e+07, 1.9095e+05, 3.9651e+06, -1.768e+07, 
    -3.5744e+06, 4.0516e+06, 2.6509e+07, 7.7394e+05, -9.5942e+06, 1.5847e+07, 
    -1.3535e+05, -1.6993e+07, -1.0447e+07, -8.4919e+06, 1.1446e+07, 
    8.7514e+06, -9.5275e+06, -1.2572e+07, -9.2076e+06, 1.0061e+07, 5.756e+05, 
    1.2177e+07, -5.9685e+06, -1.5147e+06, -3.2275e+07, 7.0358e+06, 
    -2.6773e+06, -1.6379e+07, 2.6479e+07, 2.6936e+06, 6.5404e+06, 
    -2.6148e+07, -1.0307e+06, 2.3555e+06, -1.85e+07, -1.7762e+06, 1.4634e+07, 
    -1.2984e+06, -2.387e+07, 1.0806e+07, -2.3812e+07, 6.2752e+06, 
    -6.7326e+06, 8.0616e+05, -1.3156e+07, 1.3675e+06, 2.5997e+06, 7.9784e+06, 
    -2.4837e+07, -3.9682e+06, -5.9513e+06, -6.5964e+06, -8.6886e+06, 
    2.0612e+07, 2.3089e+07, -1.1695e+06, 1.6059e+07, -3.6777e+06, 
    -1.3045e+07, -9.5734e+05, -8.129e+06, -1.997e+07, 1.6534e+07, 
    -2.1805e+07, 9.5996e+06, -1.1621e+07, 7.3753e+06, 1.2138e+07, 
    -8.6189e+05, 2.6657e+06, -1.3017e+07, -1.8527e+07, -1.0381e+07, 
    6.7068e+06, -1.8831e+07,
  -1.7819e+07, 1.7447e+07, 3.5726e+06, -5.4609e+06, 7.1626e+06, -3.0491e+07, 
    -2.4701e+06, 2.5821e+07, 1.9344e+07, 3.2381e+07, 6.1924e+06, 1.7152e+07, 
    -2.7967e+06, -2.114e+06, 4.6414e+06, -1.1747e+07, -5.5506e+06, 
    -3.0332e+07, 1.7702e+07, -1.921e+07, 1.8756e+06, 2.5573e+07, 9.3526e+06, 
    6.0739e+05, -47818, 5.9576e+06, 8.5423e+06, 7.2205e+06, -7.5801e+06, 
    -3.7723e+06, 1.5023e+06, -7.9397e+06, 1.9992e+07, 4.2831e+06, 
    -5.9141e+06, -8.5837e+06, 7.4047e+06, 7.8627e+06, -2.2368e+07, 
    3.2293e+07, -1.1279e+07, -7.747e+06, 3.4044e+07, -2.0075e+07, 1.5143e+07, 
    -1.5205e+06, 1.2398e+07, -1.1766e+06, -7.9475e+05, -87530, 4.1448e+06, 
    8.2102e+05, -2.9052e+07, 1.793e+07, 9.8946e+06, 5.017e+06, 3.4707e+06, 
    -1.7575e+06, 3.7855e+06, -3.7686e+06, -4.0855e+06, -1.9283e+07, 
    4.8644e+06, 1.0206e+07, 2.5668e+07, 5.8166e+06, -8.0716e+06, 3.3592e+07, 
    -6.9579e+05, -1.0254e+07, -1.3555e+06, -2.4528e+05, 1.103e+06, 
    4.0544e+06, -1.7913e+07, 1.4148e+07, 5.2548e+06, 2.9506e+06, 1.1744e+07, 
    1.5884e+07, 1.6334e+06, 1.9022e+06, 3.384e+06, -1.0168e+07, -9.7452e+05, 
    1.0843e+07, -9.707e+06, -7.2039e+06, 4.9833e+06, -1.9075e+05, 
    -1.1159e+07, 3.0914e+07, -6.801e+06, -1.0348e+06, -1.0293e+07, 
    2.3841e+07, 1.9053e+07, 9.0335e+06, 8.7109e+06, -2.3439e+07,
  1.506e+07, 2.5828e+06, -9.8296e+06, -3.4755e+06, 4.191e+06, -1.705e+07, 
    -1.8948e+07, -1.6505e+07, -3.0894e+07, 1.0227e+07, 2.7068e+07, 
    -2.9449e+07, 1.3577e+07, -9.6618e+06, -2.2101e+07, 5.792e+06, 1.5735e+07, 
    1.6734e+07, -1.6385e+07, 9.1774e+06, -1.8891e+06, -1.2909e+07, 
    -2.6953e+06, -2.2467e+07, 1.0284e+07, -1.758e+07, -2.3354e+07, 
    6.8472e+06, 3.4707e+07, 3.2545e+07, -8.3403e+06, 1.042e+07, -8.253e+06, 
    9.046e+06, 2.4171e+06, 2.8562e+07, -1.7818e+07, 7.6477e+05, -2.4935e+07, 
    2.3834e+06, -3.1793e+06, 1.9794e+07, 1.4359e+07, 4.5013e+06, 1.5709e+07, 
    8.5415e+06, -1.3459e+07, 2.3825e+07, 1.8259e+07, 2.383e+07, -2.9516e+07, 
    -1.4522e+07, -1.284e+07, 2.3063e+07, -4.5359e+06, 4.9899e+06, 3.1974e+07, 
    2.6115e+07, -2.8535e+07, -2.2859e+07, -2.2671e+07, -1.9045e+07, 
    -1.3244e+07, -2.5487e+07, 1.1098e+07, -1.7926e+07, 4.5231e+06, 
    2.3848e+07, 6.1116e+06, -1.8714e+07, -3.9602e+07, -1.6371e+07, 
    -1.3249e+07, -9.8563e+06, -2.7855e+07, 1.216e+07, -2.1723e+07, 
    -1.7653e+07, 6.3072e+06, -2.5786e+06, -3.8938e+07, -1.81e+07, 
    -4.0532e+06, -2.0013e+06, -4.013e+07, 3.1855e+06, -2.3098e+07, 
    1.4245e+07, 2.3669e+07, 4.9817e+06, 2.1941e+07, -6.2021e+06, -6.4214e+06, 
    -2.7225e+07, 3.972e+07, -8.0436e+06, -8.7891e+06, 1.4418e+07, 
    -7.5563e+06, -7.8953e+06 ;

 v_gns =
  1061.9, 324.61, 1011.7, 5335.5, -604.54, 491.7, -543.49, 1964.9, 1577.2, 
    -4665.8, 2975.8, 4705.6, 193.89, -1525.8, 562.53, -5440, -1116.2, 
    -341.31, -4233.5, 7326.9, 1831.9, 2372.9, 4709, 23.192, -740.2, 815.7, 
    -6526.2, 661.11, 2498.6, -1107.4, -8600, -696.78, -1807.5, 2102.2, 
    2622.9, -1443.2, 1451.8, -247.37, 481.01, -4374.2, 909.8, 4.93, -2181.1, 
    465.36, -7541.4, -1881.2, 131.59, -745.02, -1719.6, -5005.3, -104.64, 
    1813.8, -5858.1, 1198.6, 90.587, 6280.1, 1575.5, -69.658, -1742, -1236.7, 
    4296.5, -3908, 6879.7, 112.95, -75.174, 2563.9, -2308, 3045.9, -63.396, 
    2015.9, -3825.1, -128.92, 223.12, -167.23, -3437.6, 2184.1, -5706.3, 
    -7956.5, -1092.8, 3874, -2378.3, -1078.3, -2649.6, -870.65, -4784.6, 
    -56.3, 3663.5, -1718.5, 3133.3, 1056, -3937.3, -951.68, -4358.5, 7429.4, 
    3355, 2881.4, -499.05, 236.29, 348.96, -907.66,
  565.58, -452.89, -1321.4, 546.09, 8282.1, 2936.6, 1686.3, 2885.9, -1455.4, 
    -790.82, 3407.7, 7273.5, -451.3, -70.248, 1764.5, -3442, 2251.1, 947.81, 
    -3655.9, -5237.4, -1663.6, 2471.2, -1963.1, -54.323, -1080.9, 1134.3, 
    5345.2, -1753.1, -5198.1, -355.97, -4050.4, -25.731, 1098.3, -2232.3, 
    -401.13, -2275.6, -7939.3, -3410.3, 175.01, -6825.5, -507.51, -4.1344, 
    1597.7, -559.67, -693.82, -3280.8, -4305.9, -5266, -617.86, -2842.9, 
    738.05, -2352.9, -5557.8, 1214.2, 163.29, 6517.6, -1261.9, 203.92, 
    6977.9, 1490.9, -5804.2, -1020.9, 2637.4, -448.93, 1594.8, 2497.5, 
    -498.65, 151.37, -244.59, -28.891, -5429.2, 123.15, -1488.2, 773.17, 
    -861.01, -1905.9, 1723.5, -705.48, -1802.2, -4581.1, -221.6, 543.98, 
    3404, -324.58, -4413, 7384, 3082.4, -913.84, -1081.3, 1269.2, -4541.4, 
    2311.7, 2252.9, -1367, -1012.8, -42.785, -281.17, -85.491, 1620.7, 5817,
  -3276.7, 4752.8, -4296.9, -1355, 3098.4, -1510.9, -876.48, 4026.3, -2162.6, 
    -257.43, -3491.4, 696.81, -821.04, 311.49, 7285.7, -1057.5, 6223, 
    -1325.2, 3753.4, 2158.2, -4538.1, 1497.1, -6039.9, 304, -780.39, -8016.9, 
    -2041.5, 2533.5, -7395.1, -3476.8, -1224.8, 667.31, 2806.2, 5832.8, 
    -9026.8, -8337.8, -2818.8, -6421.1, -1488.3, 4460, -962.95, -147.73, 
    3163, 376.04, 2156.8, 4136.3, -5495.4, -1332.5, -1326.2, 1095.1, 944.51, 
    -2216.1, -324.55, -85.56, -2.7591, 2127, 2723, 1474.5, 1064.6, -5466, 
    276.96, -2627.7, -2242.5, -5799.3, 11.514, 1985.9, -3311.3, -4440.7, 
    2838.3, -1018.4, 975.51, -1713.9, -9296.5, 506.6, -2620, 121.72, 7167.4, 
    -1454.4, -6107.9, 814.97, 5338.7, -619.07, 1499.4, -1944.9, 4058.5, 
    -1338.5, 7862.4, 2237.1, 3723.9, 3859.6, -216.39, -7188.3, -7912.4, 
    4189.6, -5511.9, -269.93, 731.47, -445.86, 4960, -555.8 ;

 r_leo =
  -2.1531e+06, -1.8341e+06, 3.7776e+06, 6.728e+06, -4.0609e+06, -3.4721e+05, 
    -7.2717e+06, -2.0994e+06, -1.3834e+05, -3.971e+06, -4.5692e+06, 
    4.1733e+06, 6.3536e+06, 3.5726e+05, 1.9664e+06, -5.6893e+06, -4.7649e+06, 
    3.3911e+06, 69391, -4.6107e+06, -4.5391e+06, 7.7122e+06, -5.9896e+06, 
    -1.3372e+06, -9.6911e+05, -4.5238e+06, -3.0931e+06, -9.5384e+05, 
    -5.1336e+06, -6.2594e+06, -4288.3, 5.1826e+06, 3.5254e+06, -3.2272e+06, 
    -3.8268e+06, 2.3577e+06, 2.6724e+06, 1.5203e+05, 4.0518e+06, -9.0474e+06, 
    2.8871e+06, -3.5619e+06, 2.4814e+05, 86752, -2.8319e+05, -7.0723e+06, 
    -2.5784e+06, -1.9222e+06, -7.63e+06, 1.8038e+06, -2.4768e+06, 6.6213e+06, 
    -4.4075e+06, -2.5364e+06, 1.3771e+06, 3.4509e+06, -7.8239e+05, 
    -1.0503e+06, 1.3252e+06, -2.5144e+06, 2.5617e+06, -6.0616e+06, 
    -2.4339e+06, -4.9928e+06, 3.5229e+06, 5.624e+06, 6.8588e+06, -1.9757e+06, 
    9.8235e+05, -8.1745e+05, -3.5405e+06, 6.503e+06, 6.0225e+05, 1.8167e+06, 
    -4.3262e+06, -77638, -3.5476e+06, 1.3041e+06, 2.1892e+06, -2.4185e+06, 
    1.5419e+06, -3.8091e+06, 4.4264e+06, -5.6891e+06, -7.173e+05, 4.8093e+06, 
    -1.9107e+06, 3.6454e+05, -5.4895e+06, 7.601e+06, -1.255e+06, -1.0891e+06, 
    2.66e+06, 1.8613e+06, 1.6527e+06, 2.0663e+06, 1.3932e+06, 2.0045e+06, 
    7.9545e+05, -2.5773e+06,
  1.4643e+06, 4.1801e+06, 1.3637e+06, -3.2356e+06, -2.7088e+06, 5.0989e+05, 
    2.4406e+06, 4.2267e+06, -1.2544e+06, -4.7657e+06, 2.4018e+06, 
    -4.9021e+06, 2.8798e+06, 1.234e+06, -1.6052e+06, -6.1866e+06, 4.4885e+06, 
    2.4504e+06, -2.3339e+06, -2.2661e+06, 4.4025e+06, -8.3537e+05, 
    2.6194e+06, 2.7283e+06, 3.3213e+05, 5.5581e+06, -5.3128e+06, 4.2406e+06, 
    -6.2358e+06, -2.0571e+06, 7921.8, 4.8862e+06, -2.9545e+06, -1.4188e+06, 
    6.3037e+06, 3.0095e+05, -1.9374e+06, 7.8691e+05, -5.8e+06, -4.9958e+05, 
    5.4834e+06, -6.0579e+06, -4.0119e+06, -89321, -9.0577e+05, -3.2377e+06, 
    -4.4408e+05, -4.7343e+05, 1.5589e+06, -6.5228e+06, -6.8226e+06, 
    5.5554e+06, 5.4168e+06, 1.3434e+06, 4.8629e+05, -2.0079e+06, 6.971e+06, 
    6.0407e+06, 4.6574e+06, 6.9076e+06, 7.1986e+06, -2.8025e+06, -2.9621e+06, 
    4.761e+06, 7.8758e+06, 5.1879e+06, -2.3708e+06, -1.8517e+06, -5.608e+06, 
    -2.8988e+06, -5.2791e+06, 1.9144e+05, 9.5207e+06, -1.4462e+06, 
    -1.0238e+06, -3752.3, -3.9733e+06, 1.057e+05, -3.9965e+06, -4.8077e+06, 
    -8.291e+06, 2.2193e+06, 2.5102e+06, 1.3038e+06, -7.4019e+05, -9.0915e+05, 
    -2.7916e+06, 8.045e+06, -6.969e+06, 2.3431e+06, -2.6103e+06, -2.8958e+06, 
    3.3292e+06, -1.7187e+06, 8.5691e+05, -5.9008e+06, -5.0322e+06, 
    -2.4476e+06, 2.3942e+06, 7.0458e+06,
  -7.5336e+06, 8.5747e+06, -5.9266e+06, 1.2652e+06, -8.3566e+06, 7.4892e+06, 
    -6.1684e+06, 5.8128e+06, 6.7079e+06, -1.2278e+05, -5.7049e+06, 7.046e+06, 
    -3.077e+05, -6.722e+06, -8.7072e+06, 3.5882e+06, -6.3357e+06, 
    -6.7977e+06, -9.4622e+06, 7.2598e+06, 2.8181e+06, 1.8976e+06, 
    -3.9915e+06, -7.4097e+06, 6.2825e+06, -1.3887e+06, 4.19e+06, -4.8789e+06, 
    3.5273e+06, 5.3631e+06, -7.233e+06, 9.7335e+05, -5.9014e+06, -7.0007e+06, 
    -1.3738e+06, 7.4698e+06, 5.5428e+06, -6.4638e+06, -4.5127e+06, 
    -2.6681e+05, -3.0104e+06, -1.7356e+06, -7.7523e+06, -6.3383e+06, 
    -9.4108e+06, -2.1142e+06, 8.1869e+06, -8.8532e+06, -4.8771e+05, 
    6.2121e+06, -3.4777e+06, -1.311e+06, 2.825e+06, -7.9736e+06, 6.6603e+06, 
    4.98e+06, -1.1598e+06, -2.5658e+06, -5.4949e+06, 1.8535e+06, -3.7273e+05, 
    -3.212e+06, 4.9773e+06, 4.1612e+06, 4.1805e+06, -4.3339e+06, 6.0086e+06, 
    9.2733e+06, -6.249e+06, -8.3923e+06, -4.3808e+06, -2.409e+06, 
    -1.0039e+06, 7.2752e+06, -5.2878e+06, -7.5873e+06, 7.022e+06, 
    -9.7217e+06, -5.9016e+06, -6.7664e+06, -1.3966e+06, 7.5042e+06, 
    -4.0381e+06, 5.8764e+06, 8.823e+06, -5.286e+06, 8.0868e+06, 5.747e+06, 
    2.3232e+06, 3.89e+06, 8.9857e+06, 6.6141e+06, 4.7481e+06, 9.1232e+06, 
    -6.257e+06, -2.4113e+06, 3.9649e+06, -8.3938e+06, 8.9565e+06, 3.4416e+05 ;

 v_leo =
  3154.2, 1401.1, 30.745, -304.67, -253, -2766.8, 217.04, -1695.1, -422.28, 
    -1758.6, 6204.7, -1131.6, -868.08, 264.84, 306.55, 4192.7, 1187.8, 
    1693.5, -653.51, -4330.1, 127.09, -2116.2, 1460.2, 20.614, 4957.9, 
    -415.89, -639.43, 5155.8, -795.55, 2686.3, 1406.7, 3967.6, -2583.3, 
    1397.7, -5142.6, 1072.5, -332.28, -1456.3, -1156.6, -2746.8, -1011.4, 
    -2675.3, 377.96, 1289.8, 1822.1, -1260.8, -2438.5, 283.24, 2217.2, 
    -1.5899, -254.46, 13.687, 1042, 6600.6, -2419.1, 2170.5, 445.01, 4763.2, 
    -230, -148.26, -327.11, -2428.1, 404.21, 207.07, -2084.2, -21.335, 
    -4454.1, 3311.5, 5427.6, 569.96, -111.94, 149.61, 587.91, 280.56, 582.88, 
    2211.8, -290.24, 15.019, 5497.8, -315.56, 13.126, 2157.6, 1010.7, -1303, 
    35.969, -2560.4, 181.7, -3338.9, 59.833, 4177, -2570.1, -2373.9, -2716.8, 
    47.782, -2729.8, -1349.2, 1394.2, -1711.6, 2315.2, -1763.7,
  3583.4, 167.92, 480.03, -1728.8, -5475.1, 478.25, -280.29, 2072, 1708.6, 
    -4119.3, -3562.9, 902.61, 4750.9, -63.31, 228.45, 578.25, 2931.7, 
    -4595.9, -883.5, -3495.5, 268.79, -37.156, 3544.4, -37.984, 7972.5, 
    183.93, 477.75, -3448.6, 1487.9, 2619.1, 514.16, -4608.8, -804.81, 
    580.72, 1529.1, 6272.1, 403.74, 763.05, -757.24, -3261.6, 3729.2, 
    -661.62, -3523.6, -2758.7, 6140.9, -7632.1, -1103.3, -848.28, 688.12, 
    9.3916, -788.87, -88.834, 1626.9, -1037.4, 1634.5, 5994.7, 258.35, 
    898.47, -364.82, -163.11, 87.65, 866.06, 576.86, -463.34, 4732.3, 
    -356.69, 3528.3, 2891.1, -7000.7, -492.28, 88.989, -480.15, 1631.9, 
    -127.24, -1003.6, -3268.4, -259.04, 248.19, -1226.3, -4484.8, 73.837, 
    844.75, -192.15, 744.27, 21.48, -156.99, 515.58, 6127.4, -848.74, 
    -5010.4, 1509.3, -2493.6, 2216.4, -46.612, -6716, 1588, 677.56, 2028.8, 
    -1514.1, -397.57,
  -5417.8, 5050.3, 2285.6, -2861.9, 824.34, -2006.5, -253.46, 1886.8, 984.93, 
    3941.6, 5895.9, 1012.7, -7918.8, -2529.1, 639.23, -4861.9, -7886.8, 
    -4420.4, 3151.6, -1595.3, 4578, 2875.3, 1906, 336.2, -112.35, 2214.7, 
    780.56, 3670.3, -8217.6, -8723.4, 268.72, -891.14, 2603.1, 7103.2, 
    -968.48, -6464.3, 2509, 4918.4, -2003.6, 3012.7, -1892.6, -7757.6, 
    5086.5, -4747.2, 3434.6, -5342.9, 1122.7, -9160.7, -9420.9, -7024.4, 226, 
    599.68, -3307.2, 2049.4, 2231, 2163.6, 7787.4, -8462.2, 239.59, -2186.4, 
    -516.5, -1279.9, 917.05, 2477.8, 3433.5, 2968.7, -2779.9, 5364.5, 
    -3294.1, -2191.5, -58.862, -23.672, 119.33, 3799.3, -1445.8, 5941.4, 
    1112.7, 1505.4, 1492.1, 1397.2, 145.94, 136.75, 2637.4, -4366, -99.884, 
    5129.2, -2375.1, -1454.1, 7542.1, -64.802, -7406.7, 2718.1, -915.3, 
    -142.47, -5611.2, 3511.9, 3669.3, 7093.8, 1361.4, -3771.7 ;

 phase_qual =
  46.848, 74.886, 19.119, 2.2919, 50.294, 82.231, 35.128, 70.113, 87.322, 
    76.116, 58.678, 77.308, 21.025, 20.803, 44.893, 19.02, 31.159, 77.667, 
    72.413, 84.786, 22.888, 63.943, 15.858, 44.551, 11.619, 46.159, 50.729, 
    12.26, 90.983, 72.711, 8.6772, 63.504, 41.963, 20.827, 29.584, 64.197, 
    53.021, 18.743, 77.057, 76.478, 22.896, 46.45, 89.209, 44.401, 48.442, 
    6.7794, 42.881, 49.971, 32.987, 92.172, 66.371, 23.341, 80.265, 90.292, 
    13.622, 9.3361, 95.788, 54.332, 61.635, 63.717, 45.937, 66.85, 21.654, 
    82.013, 64.62, 65.672, 13.532, 96.585, 0.0099449, 51.274, 90.894, 28.201, 
    25.286, 56.595, 73.789, 36.363, 46.475, 37.216, 49.856, 59.629, 89.103, 
    49.109, 0.63777, 28.424, 92.265, 20.981, 70.217, 45.605, 71.646, 12.546, 
    57.121, 71.143, 24.793, 57.225, 94.888, 60.134, 59.215, 37.313, 19.402, 
    67.624 ;

 lat_tp =
  18.184, -25.924, -34.216, 65.838, 63.081, -38.987, 54.453, -49.596, 12.452, 
    -69.343, 74.07, -42.571, -50.826, -34.638, 84.534, 20.465, 36.506, 
    16.846, -82.772, -35.584, 83.277, -10.314, -85.85, 41.812, -75.737, 
    79.321, -77.406, 69.441, -78.997, -10.755, 0.91548, 51.884, 36.137, 
    67.782, 76.011, 70.268, -39.813, -12.38, -64.822, -60.162, -46.162, 
    47.964, -55.85, -43.652, 77.38, -82.985, 35.178, -2.1015, -44.967, 
    -16.177, 66.877, 0.06429, -76.737, -88.916, 12.595, 25.103, -34.806, 
    25.54, -34.793, 64.79, 49.416, 25.727, 57.185, 21.283, 18.549, -52.302, 
    31.132, 35.968, -86.425, 7.5904, 35.723, 72.109, 82.23, 23.848, -78.115, 
    -45.278, 60.385, 53.778, -59.377, 54.502, -70.832, -2.309, -65.839, 
    79.762, 1.7363, -65.176, 43.892, -35.08, -18.509, 80.422, -18.126, 
    -76.81, -50.816, 65.119, 78.253, 10.372, 67.637, 13.206, 9.1135, 34.158 ;

 lon_tp =
  61.38, 67.235, 112.93, -40.659, -54.702, -172.08, 100.06, 128.21, 55.448, 
    164.89, -11.394, -48.575, 59.856, 115.6, -117.41, 44.734, 0.82563, 
    -55.544, -12.997, 41.815, -162.55, 62.081, -158.66, 125.75, -95.707, 
    10.455, 85.003, -147.68, 104.88, 83.423, 46.731, -81.76, 74.651, 15.847, 
    -155.22, -30.186, -116.7, 107.06, 47.017, -168.24, 129.21, 14.995, 
    141.81, 163.49, 17.244, 25.056, 87.275, 67.104, -43.276, -117.67, 
    -11.981, -67.62, 81.434, 137.98, -171.71, 55.519, -125.84, 20.647, 
    93.409, -105.43, 125.3, -90.8, 129.15, -57.514, 43.744, 31.168, -98.598, 
    129.39, 160.2, -132.34, -12.929, -117.89, -2.1006, 105.38, 87.862, 
    -74.88, -74.097, -54.904, -28.855, -6.1142, -121.38, -138.35, -52.416, 
    -177.92, 53.287, 124.66, -3.0822, -88.273, -12.076, -155.92, -63.348, 
    -48.51, 101.13, -79.69, 165.39, 113.42, -123.32, -33.73, -80.103, 122.75 ;

 azimuth_tp =
  42.091, 210.89, 171.94, 117.34, 236.33, 91.16, 311.42, 229.68, 69.031, 
    57.041, 216.56, 139.01, 245.86, 15.374, 271.04, 149.68, 298.55, 124.75, 
    147.96, 267.93, 203.68, 232.15, 233.72, 265.57, 106.94, 117.69, 115.34, 
    107.16, 151.94, 133.66, 332.78, 303.84, 160.14, 302.39, 174.34, 303.39, 
    349.71, 225.3, 119.38, 120.46, 89.099, 329.59, 198.34, 328.84, 183.7, 
    89.333, 27.49, 84.359, 289.73, 57.023, 147.54, 54.197, 287.04, 179.5, 
    280.13, 128.96, 21.341, 246.18, 49.951, 85.947, 125.37, 351.68, 284.61, 
    219.93, 93.827, 78.854, 142.54, 321.42, 131.64, 18.876, 298.64, 98.321, 
    44.255, 240.81, 234.6, 42.466, 307.24, 210.24, 23.972, 288.29, 89.038, 
    64.474, 171.51, 149.77, 187.57, 261.32, 174.39, 298.65, 26.911, 90.04, 
    197.05, 14.716, 294.04, 156.72, 11.249, 324.1, 106.5, 126.17, 173.53, 
    138.04 ;

 impact_L1 =
  6.3467e+06, 6.2341e+06, 6.5652e+06, 6.2906e+06, 6.5913e+06, 6.2454e+06, 
    6.5777e+06, 6.3437e+06, 6.3211e+06, 6.3052e+06, 6.3051e+06, 6.3361e+06, 
    6.2147e+06, 6.2087e+06, 6.4019e+06, 6.2984e+06, 6.4401e+06, 6.3955e+06, 
    6.5033e+06, 6.514e+06, 6.479e+06, 6.5176e+06, 6.385e+06, 6.4863e+06, 
    6.3568e+06, 6.4958e+06, 6.3616e+06, 6.2893e+06, 6.5892e+06, 6.4833e+06, 
    6.3338e+06, 6.3298e+06, 6.5306e+06, 6.3128e+06, 6.2847e+06, 6.3709e+06, 
    6.5594e+06, 6.3351e+06, 6.4386e+06, 6.4357e+06, 6.4975e+06, 6.5191e+06, 
    6.3052e+06, 6.5181e+06, 6.3901e+06, 6.4102e+06, 6.2822e+06, 6.2355e+06, 
    6.4258e+06, 6.511e+06, 6.2994e+06, 6.5351e+06, 6.5375e+06, 6.5002e+06, 
    6.5354e+06, 6.5068e+06, 6.3952e+06, 6.403e+06, 6.2061e+06, 6.3516e+06, 
    6.297e+06, 6.3482e+06, 6.2977e+06, 6.574e+06, 6.4861e+06, 6.441e+06, 
    6.2218e+06, 6.5451e+06, 6.4598e+06, 6.5206e+06, 6.4913e+06, 6.5508e+06, 
    6.2906e+06, 6.5655e+06, 6.3361e+06, 6.2106e+06, 6.2109e+06, 6.3474e+06, 
    6.4169e+06, 6.4921e+06, 6.5781e+06, 6.5122e+06, 6.2036e+06, 6.2205e+06, 
    6.2152e+06, 6.3715e+06, 6.3696e+06, 6.5027e+06, 6.3114e+06, 6.3985e+06, 
    6.5179e+06, 6.4985e+06, 6.4898e+06, 6.5846e+06, 6.5841e+06, 6.2175e+06, 
    6.3281e+06, 6.5675e+06, 6.2202e+06, 6.5426e+06 ;

 impact_L2 =
  6.5663e+06, 6.4813e+06, 6.3952e+06, 6.3995e+06, 6.5205e+06, 6.5063e+06, 
    6.3082e+06, 6.482e+06, 6.2627e+06, 6.4103e+06, 6.5729e+06, 6.4036e+06, 
    6.4244e+06, 6.2748e+06, 6.3551e+06, 6.3205e+06, 6.3807e+06, 6.333e+06, 
    6.4249e+06, 6.4022e+06, 6.2895e+06, 6.4043e+06, 6.3873e+06, 6.2077e+06, 
    6.3615e+06, 6.5845e+06, 6.2447e+06, 6.3951e+06, 6.5523e+06, 6.452e+06, 
    6.5787e+06, 6.4155e+06, 6.2804e+06, 6.3474e+06, 6.2801e+06, 6.4361e+06, 
    6.2518e+06, 6.5273e+06, 6.293e+06, 6.2664e+06, 6.4221e+06, 6.5469e+06, 
    6.4858e+06, 6.2583e+06, 6.4781e+06, 6.3014e+06, 6.3996e+06, 6.4525e+06, 
    6.5732e+06, 6.5011e+06, 6.3938e+06, 6.4578e+06, 6.2997e+06, 6.3981e+06, 
    6.2423e+06, 6.4656e+06, 6.2046e+06, 6.36e+06, 6.3492e+06, 6.5266e+06, 
    6.4921e+06, 6.3368e+06, 6.3282e+06, 6.5354e+06, 6.3068e+06, 6.3931e+06, 
    6.4504e+06, 6.238e+06, 6.4184e+06, 6.4442e+06, 6.2514e+06, 6.4487e+06, 
    6.2533e+06, 6.2491e+06, 6.2616e+06, 6.2737e+06, 6.3327e+06, 6.3742e+06, 
    6.4625e+06, 6.2077e+06, 6.3192e+06, 6.3386e+06, 6.2809e+06, 6.2336e+06, 
    6.2922e+06, 6.2553e+06, 6.4058e+06, 6.3916e+06, 6.3456e+06, 6.247e+06, 
    6.4199e+06, 6.4268e+06, 6.2216e+06, 6.3074e+06, 6.4566e+06, 6.5404e+06, 
    6.3893e+06, 6.3286e+06, 6.2725e+06, 6.4777e+06 ;

 impact =
  6.4143e+06, 6.3427e+06, 6.3882e+06, 6.3012e+06, 6.4999e+06, 6.5327e+06, 
    6.4639e+06, 6.4916e+06, 6.4672e+06, 6.4098e+06, 6.2324e+06, 6.4234e+06, 
    6.3786e+06, 6.3119e+06, 6.441e+06, 6.2186e+06, 6.2479e+06, 6.4236e+06, 
    6.3218e+06, 6.2671e+06, 6.3487e+06, 6.5046e+06, 6.4331e+06, 6.2179e+06, 
    6.447e+06, 6.5288e+06, 6.324e+06, 6.5259e+06, 6.4146e+06, 6.4711e+06, 
    6.3549e+06, 6.2463e+06, 6.3283e+06, 6.3388e+06, 6.5377e+06, 6.4315e+06, 
    6.218e+06, 6.3561e+06, 6.3573e+06, 6.4439e+06, 6.2511e+06, 6.4866e+06, 
    6.2738e+06, 6.4121e+06, 6.3416e+06, 6.3461e+06, 6.2775e+06, 6.492e+06, 
    6.4921e+06, 6.5592e+06, 6.3831e+06, 6.4449e+06, 6.544e+06, 6.5011e+06, 
    6.5455e+06, 6.4014e+06, 6.3027e+06, 6.3472e+06, 6.3228e+06, 6.3499e+06, 
    6.5162e+06, 6.2029e+06, 6.446e+06, 6.3354e+06, 6.312e+06, 6.265e+06, 
    6.3592e+06, 6.3727e+06, 6.2739e+06, 6.2485e+06, 6.3176e+06, 6.3694e+06, 
    6.3664e+06, 6.2638e+06, 6.2075e+06, 6.529e+06, 6.4762e+06, 6.3186e+06, 
    6.518e+06, 6.277e+06, 6.2713e+06, 6.5112e+06, 6.5775e+06, 6.4266e+06, 
    6.3181e+06, 6.4906e+06, 6.2312e+06, 6.5835e+06, 6.4705e+06, 6.3644e+06, 
    6.5833e+06, 6.4787e+06, 6.2678e+06, 6.2873e+06, 6.475e+06, 6.5265e+06, 
    6.5472e+06, 6.5224e+06, 6.3858e+06, 6.3613e+06 ;

 impact_opt =
  6.4156e+06, 6.4098e+06, 6.3775e+06, 6.3284e+06, 6.4673e+06, 6.439e+06, 
    6.4496e+06, 6.5618e+06, 6.2605e+06, 6.2762e+06, 6.3376e+06, 6.499e+06, 
    6.5428e+06, 6.571e+06, 6.3498e+06, 6.4703e+06, 6.4534e+06, 6.3052e+06, 
    6.4651e+06, 6.3444e+06, 6.5104e+06, 6.5e+06, 6.32e+06, 6.3234e+06, 
    6.2302e+06, 6.4084e+06, 6.315e+06, 6.5172e+06, 6.565e+06, 6.4303e+06, 
    6.4093e+06, 6.3693e+06, 6.4391e+06, 6.3181e+06, 6.2937e+06, 6.4792e+06, 
    6.398e+06, 6.2765e+06, 6.5367e+06, 6.2993e+06, 6.4124e+06, 6.2964e+06, 
    6.2104e+06, 6.3656e+06, 6.5183e+06, 6.2055e+06, 6.3865e+06, 6.4659e+06, 
    6.5831e+06, 6.3012e+06, 6.3388e+06, 6.2708e+06, 6.5506e+06, 6.3966e+06, 
    6.4382e+06, 6.2305e+06, 6.304e+06, 6.5247e+06, 6.4773e+06, 6.2336e+06, 
    6.3723e+06, 6.3557e+06, 6.5558e+06, 6.2526e+06, 6.4141e+06, 6.2599e+06, 
    6.249e+06, 6.2246e+06, 6.2349e+06, 6.4344e+06, 6.5742e+06, 6.4847e+06, 
    6.3963e+06, 6.2626e+06, 6.4148e+06, 6.3772e+06, 6.5297e+06, 6.258e+06, 
    6.4611e+06, 6.5322e+06, 6.4379e+06, 6.3752e+06, 6.367e+06, 6.3868e+06, 
    6.2923e+06, 6.2913e+06, 6.2267e+06, 6.4585e+06, 6.4674e+06, 6.2693e+06, 
    6.5625e+06, 6.4859e+06, 6.2222e+06, 6.5578e+06, 6.3046e+06, 6.2747e+06, 
    6.429e+06, 6.3184e+06, 6.3714e+06, 6.3197e+06 ;

 bangle_L1 =
  0.047544, 0.097615, 0.087559, 0.075333, 0.09107, 0.0033325, 0.066036, 
    0.032596, 2.4718e-05, 0.035244, 0.032477, 0.01681, 0.031999, 0.023942, 
    0.022785, 0.039151, 0.015515, 0.0010231, 0.055641, 0.083262, 0.0041524, 
    0.0027358, 0.062049, 0.013235, 0.066762, 0.020452, 0.090433, 0.012671, 
    0.054819, 0.024612, 0.025625, 0.033454, 0.083472, 0.061375, 0.024976, 
    0.046941, 0.036685, 0.034274, 0.084944, 0.078026, 0.068033, 0.041151, 
    0.013411, 0.091887, 0.096848, 0.088175, 0.025899, 0.064467, 0.0071828, 
    0.018651, 0.047486, 0.074195, 0.016799, 0.032737, 0.050738, 0.071302, 
    0.06944, 0.006108, 0.076052, 0.0082807, 0.0053619, 0.063903, 0.095544, 
    0.088232, 0.0789, 0.043171, 0.052112, 0.050356, 0.03941, 0.018837, 
    0.094075, 0.043855, 0.059727, 0.021235, 0.090272, 0.021248, 0.042121, 
    0.071962, 0.088141, 0.057636, 0.06615, 0.088555, 0.053214, 0.030872, 
    0.004237, 0.011698, 0.06262, 0.083769, 0.093352, 0.027536, 0.043039, 
    0.051414, 0.034554, 0.064321, 0.075862, 0.0070635, 0.075092, 0.041979, 
    0.056163, 0.082355 ;

 bangle_L2 =
  0.08126, 0.056385, 0.091988, 0.028994, 0.00012125, 0.0050322, 0.047432, 
    0.034707, 0.065765, 0.065207, 0.040004, 0.093475, 0.08563, 0.0082613, 
    0.016305, 0.086173, 0.08004, 0.015318, 0.04271, 0.024958, 0.051163, 
    0.029557, 0.095921, 0.049454, 0.094209, 0.015285, 0.036139, 0.0078812, 
    0.0084967, 0.0066131, 0.008298, 0.018941, 0.050603, 0.018063, 0.085167, 
    0.062194, 0.049713, 0.082718, 0.075475, 0.00461, -0.00068496, 0.088179, 
    0.087278, 0.015323, 0.086152, 0.0037044, 0.062717, 0.012441, 0.022509, 
    0.058699, 0.047085, 0.028279, 0.074449, 0.061843, 0.026052, 0.016342, 
    0.070701, 0.0051497, 0.070994, 0.062166, 0.07552, 0.060585, 0.029161, 
    0.037179, 0.022066, 0.039078, 0.051859, 0.0064769, 0.069983, 0.023665, 
    0.09373, 0.070897, 0.07718, 0.073255, 0.030034, 0.0056779, 0.047966, 
    0.037851, 0.069977, 0.040802, -0.00041461, 0.063488, 0.043278, 0.037636, 
    0.093012, 0.053188, 0.077202, 0.052399, 0.012986, 0.063536, 0.089623, 
    0.014637, 0.043381, 0.010652, 0.073737, 0.029499, 0.0068787, 0.060431, 
    0.059266, 0.027051 ;

 bangle =
  0.0026314, 0.085925, 0.075215, 0.0094704, 0.062516, 0.012931, 0.015797, 
    0.0025448, 0.037404, 0.047348, 0.095404, 0.092432, 0.034815, 0.055743, 
    0.021134, 0.029665, 0.052632, 0.034162, 0.00295, 0.096904, 0.079807, 
    0.024642, 0.079431, 0.048675, 0.014292, 0.059755, 0.083655, 0.034585, 
    0.055431, 0.052164, 0.034183, 0.072851, 0.030543, 0.084519, 0.058147, 
    0.027461, 0.0071483, 0.011612, 0.039055, 0.043856, 0.03256, 0.059944, 
    0.061532, 0.053259, 0.035061, 0.024432, 0.060386, 0.0281, 0.090899, 
    0.091214, 0.037614, 0.0081933, 0.034482, 0.021594, 0.012244, 0.013376, 
    0.0011179, 0.06694, 0.020318, 0.059523, 0.079821, 0.034193, 0.053369, 
    0.087447, 0.06789, 0.012138, 0.061246, 0.06113, 0.034773, 0.011066, 
    0.084047, 0.067892, 0.05531, 0.090125, 0.081876, 0.00065058, 0.040538, 
    0.020777, 0.018736, 0.026213, 0.087347, 0.013739, 0.055633, 0.054137, 
    0.055261, 0.082622, 0.0474, 0.01994, 0.066653, 0.0054888, 0.094699, 
    0.093515, 0.049462, 0.071713, 0.006026, 0.045837, 0.053513, 0.024679, 
    0.029185, 0.048491 ;

 bangle_opt =
  0.059703, 0.034954, 0.030301, 0.086443, 0.084895, 0.027624, 0.080054, 
    0.021671, 0.056487, 0.010591, 0.091062, 0.025613, 0.020981, 0.030064, 
    0.096933, 0.060983, 0.069984, 0.058952, 0.0030557, 0.029533, 0.096228, 
    0.043712, 0.0013287, 0.072961, 0.0070031, 0.094008, 0.0060664, 0.088464, 
    0.0051736, 0.043465, 0.050014, 0.078613, 0.069777, 0.087533, 0.092151, 
    0.088928, 0.02716, 0.042553, 0.013127, 0.015743, 0.023598, 0.076413, 
    0.018162, 0.025006, 0.092919, 0.0029363, 0.069239, 0.048321, 0.024269, 
    0.040423, 0.087026, 0.049536, 0.0064421, -0.00039186, 0.056567, 0.063586, 
    0.02997, 0.06383, 0.029977, 0.085854, 0.077228, 0.063936, 0.081587, 
    0.061442, 0.059908, 0.020153, 0.066969, 0.069682, 0.0010059, 0.053759, 
    0.069544, 0.089961, 0.09564, 0.062882, 0.0056687, 0.024094, 0.083383, 
    0.079675, 0.016183, 0.080082, 0.0097554, 0.048204, 0.012557, 0.094256, 
    0.050474, 0.012929, 0.074128, 0.029816, 0.039114, 0.094626, 0.039329, 
    0.0064008, 0.020987, 0.086039, 0.093408, 0.05532, 0.087452, 0.05691, 
    0.054614, 0.068667 ;

 bangle_L1_sigma =
  0.0063597, 0.006514, 0.0077178, 0.0036712, 0.0033012, 0.00020866, 
    0.0073788, 0.0081204, 0.0062034, 0.009087, 0.0044423, 0.0034627, 
    0.0063195, 0.0077884, 0.001649, 0.0059211, 0.0047643, 0.0032791, 
    0.0044001, 0.0058442, 0.00045988, 0.0063782, 0.00056213, 0.0080558, 
    0.0022209, 0.005018, 0.0069821, 0.0008516, 0.0075058, 0.0069405, 
    0.0059737, 0.0025884, 0.0067093, 0.00516, 0.0006529, 0.0039472, 
    0.0016679, 0.0075631, 0.0059813, 0.00030977, 0.0081469, 0.0051376, 
    0.0084788, 0.0090501, 0.0051968, 0.0054027, 0.0070419, 0.0065105, 
    0.0036023, 0.0016422, 0.0044268, 0.0029609, 0.0068881, 0.0083778, 
    0.0002184, 0.0062053, 0.001427, 0.0052865, 0.0072036, 0.0019646, 
    0.0080437, 0.0023502, 0.0081452, 0.0032272, 0.005895, 0.0055637, 
    0.0021447, 0.0081517, 0.0089633, 0.0012557, 0.0044019, 0.0016364, 
    0.0046872, 0.0075189, 0.0070574, 0.0027696, 0.0027903, 0.0032959, 
    0.0039822, 0.0045814, 0.0015445, 0.0010973, 0.0033615, 5.4718e-05, 
    0.0061465, 0.008027, 0.0046613, 0.0024168, 0.0044243, 0.00063437, 
    0.0030735, 0.0034644, 0.0074071, 0.0026429, 0.0091002, 0.0077308, 
    0.0014934, 0.0038538, 0.002632, 0.0079766 ;

 bangle_L2_sigma =
  0.001109, 0.0055563, 0.0045301, 0.0030915, 0.0062268, 0.0024018, 0.008205, 
    0.0060515, 0.0018188, 0.0015029, 0.0057058, 0.0036624, 0.0064777, 
    0.00040507, 0.0071411, 0.0039436, 0.0078661, 0.0032869, 0.0038982, 
    0.0070593, 0.0053664, 0.0061164, 0.0061578, 0.006997, 0.0028177, 
    0.0031009, 0.0030388, 0.0028233, 0.0040033, 0.0035217, 0.0087678, 
    0.0080055, 0.0042194, 0.0079672, 0.0045934, 0.0079934, 0.0092139, 
    0.0059361, 0.0031453, 0.0031739, 0.0023475, 0.0086837, 0.0052257, 
    0.0086641, 0.0048399, 0.0023537, 0.00072428, 0.0022226, 0.0076336, 
    0.0015024, 0.0038873, 0.0014279, 0.0075628, 0.0047292, 0.0073807, 
    0.0033979, 0.00056228, 0.0064862, 0.0013161, 0.0022645, 0.0033032, 
    0.0092658, 0.0074988, 0.0057946, 0.0024721, 0.0020776, 0.0037556, 
    0.0084684, 0.0034683, 0.00049732, 0.0078683, 0.0025905, 0.001166, 
    0.0063447, 0.006181, 0.0011189, 0.0080948, 0.0055392, 0.0006316, 
    0.0075956, 0.0023459, 0.0016987, 0.0045188, 0.0039459, 0.0049419, 
    0.0068851, 0.0045946, 0.0078687, 0.00070903, 0.0023723, 0.0051918, 
    0.00038772, 0.0077472, 0.0041291, 0.00029637, 0.0085392, 0.0028059, 
    0.0033241, 0.004572, 0.003637 ;

 bangle_sigma =
  0.0034782, 0.00080743, 0.00866, 0.0021487, 0.0092783, 0.0010771, 0.0089561, 
    0.0034083, 0.002872, 0.0024943, 0.0024914, 0.003227, 0.00034878, 
    0.00020609, 0.0047883, 0.0023334, 0.0056934, 0.0046352, 0.0071927, 
    0.0074464, 0.0066155, 0.0075312, 0.0043871, 0.0067878, 0.0037188, 
    0.0070134, 0.0038329, 0.0021167, 0.0092288, 0.0067169, 0.003172, 
    0.0030774, 0.007839, 0.0026755, 0.0020082, 0.0040525, 0.0085213, 
    0.0032025, 0.0056584, 0.005589, 0.0070538, 0.0075669, 0.0024938, 
    0.0075424, 0.0045081, 0.0049839, 0.0019484, 0.00084195, 0.0053535, 
    0.007374, 0.0023579, 0.0079471, 0.0080037, 0.0071178, 0.0079526, 
    0.0072756, 0.0046291, 0.0048148, 0.00014537, 0.0035957, 0.0022996, 
    0.0035148, 0.002316, 0.0088681, 0.0067844, 0.0057156, 0.00051682, 
    0.008182, 0.0061613, 0.0076033, 0.006907, 0.0083194, 0.0021483, 
    0.0086666, 0.0032278, 0.0002503, 0.00025788, 0.0034963, 0.0051421, 
    0.0069268, 0.008966, 0.0074026, 8.6093e-05, 0.00048688, 0.00036065, 
    0.0040678, 0.0040209, 0.0071785, 0.0026422, 0.0047064, 0.0075388, 
    0.0070782, 0.0068711, 0.0091188, 0.0091087, 0.00041388, 0.0030385, 
    0.0087142, 0.00047863, 0.0081232 ;

 bangle_opt_sigma =
  0.0091566, 0.0070321, 0.0048801, 0.0049866, 0.0080132, 0.0076585, 0.002705, 
    0.007051, 0.0015682, 0.0052569, 0.0093226, 0.0050894, 0.0056095, 
    0.001871, 0.0038781, 0.0030124, 0.0045184, 0.0033252, 0.0056214, 
    0.0050541, 0.0022378, 0.0051069, 0.0046824, 0.00019183, 0.0040379, 
    0.0096137, 0.001118, 0.0048787, 0.0088084, 0.0062991, 0.0094687, 
    0.0053864, 0.0020108, 0.0036859, 0.0020037, 0.005903, 0.0012941, 
    0.0081831, 0.0023239, 0.0016608, 0.0055529, 0.0086736, 0.0071438, 
    0.0014572, 0.0069537, 0.0025347, 0.0049888, 0.0063133, 0.0093302, 
    0.0075263, 0.0048461, 0.0064456, 0.0024916, 0.0049516, 0.0010578, 
    0.0066412, 0.00011615, 0.0039991, 0.0037305, 0.0081642, 0.0073015, 
    0.0034192, 0.0032038, 0.0083851, 0.0026696, 0.0048281, 0.0062595, 
    0.00094927, 0.005459, 0.006106, 0.0012858, 0.0062181, 0.0013317, 
    0.0012269, 0.0015405, 0.0018425, 0.0033171, 0.0043555, 0.0065636, 
    0.00019319, 0.0029807, 0.0034644, 0.0020229, 0.00084053, 0.0023052, 
    0.0013834, 0.0051458, 0.0047899, 0.0036407, 0.0011742, 0.0054985, 
    0.0056696, 0.00054109, 0.0026855, 0.0064156, 0.0085107, 0.0047322, 
    0.0032157, 0.0018119, 0.0069432 ;

 bangle_L1_qual =
  53.583, 35.666, 47.039, 25.312, 74.972, 83.176, 65.972, 72.905, 66.795, 
    52.438, 8.0904, 55.849, 44.642, 27.975, 60.262, 4.6453, 11.973, 55.893, 
    30.458, 16.768, 37.165, 76.156, 58.276, 4.4642, 61.752, 82.199, 30.995, 
    81.465, 53.66, 67.769, 38.714, 11.576, 32.084, 34.7, 84.434, 57.887, 
    4.5093, 39.031, 39.313, 60.978, 12.773, 71.66, 18.456, 53.026, 35.404, 
    36.527, 19.365, 73.004, 73.016, 89.796, 45.772, 61.237, 86.01, 75.28, 
    86.363, 50.342, 25.675, 36.796, 30.708, 37.48, 79.051, 0.73518, 61.506, 
    33.858, 27.996, 16.254, 39.789, 43.174, 18.473, 12.128, 29.412, 42.341, 
    41.591, 15.944, 1.876, 82.243, 69.048, 29.638, 79.494, 19.258, 17.816, 
    77.799, 94.38, 56.659, 29.527, 72.661, 7.8109, 95.868, 67.63, 41.094, 
    95.834, 69.685, 16.945, 21.83, 68.748, 81.619, 86.793, 80.608, 46.443, 
    40.33 ;

 bangle_L2_qual =
  53.904, 52.446, 44.372, 32.104, 66.828, 59.741, 62.406, 90.443, 15.124, 
    19.046, 34.41, 74.76, 85.709, 92.753, 37.45, 67.566, 63.358, 26.298, 
    66.283, 36.105, 77.588, 74.993, 30.001, 30.861, 7.5601, 52.088, 28.753, 
    79.303, 91.261, 57.575, 52.321, 42.329, 59.78, 29.536, 23.426, 69.806, 
    49.503, 19.136, 84.184, 24.837, 53.094, 24.107, 2.6035, 41.392, 79.57, 
    1.3874, 46.629, 66.484, 95.765, 25.296, 34.698, 17.712, 87.647, 49.148, 
    59.541, 7.6219, 26.006, 81.179, 69.316, 8.3878, 43.077, 38.92, 88.961, 
    13.161, 53.518, 14.984, 12.248, 6.147, 8.7219, 58.608, 93.559, 71.18, 
    49.087, 15.654, 53.697, 44.289, 82.418, 14.509, 65.279, 83.054, 59.474, 
    43.803, 41.751, 46.703, 23.079, 22.831, 6.6649, 64.613, 66.858, 17.328, 
    90.623, 71.486, 5.5545, 89.439, 26.155, 18.672, 57.253, 29.607, 42.852, 
    29.92 ;

 bangle_qual =
  48.063, 97.639, 87.682, 75.577, 91.158, 4.2896, 66.373, 33.264, 1.0146, 
    35.885, 33.145, 17.633, 32.673, 24.695, 23.549, 39.754, 16.352, 2.0031, 
    56.08, 83.428, 5.1014, 3.6988, 62.424, 14.094, 67.091, 21.239, 90.527, 
    13.536, 55.267, 25.358, 26.362, 34.113, 83.635, 61.757, 25.719, 47.466, 
    37.311, 34.925, 85.093, 78.244, 68.349, 41.733, 14.268, 91.967, 96.879, 
    88.292, 26.632, 64.819, 8.1018, 19.456, 48.006, 74.45, 17.623, 33.403, 
    51.226, 71.586, 69.743, 7.0376, 76.289, 9.1888, 6.2989, 64.26, 95.588, 
    88.348, 79.109, 43.733, 52.586, 50.847, 40.01, 19.64, 94.134, 44.411, 
    60.125, 22.015, 90.368, 22.028, 42.694, 72.239, 88.258, 58.056, 66.485, 
    88.669, 53.677, 31.556, 5.1851, 12.572, 62.99, 83.93, 93.418, 28.254, 
    43.603, 51.895, 35.202, 64.674, 76.101, 7.9836, 75.339, 42.553, 56.597, 
    82.53 ;

 bangle_opt_qual =
  81.445, 56.817, 92.067, 29.697, 1.1102, 5.9725, 47.953, 35.354, 66.104, 
    65.552, 40.598, 93.539, 85.772, 9.1696, 17.133, 86.309, 80.238, 16.157, 
    43.277, 25.701, 51.647, 30.255, 95.962, 49.955, 94.266, 16.124, 36.771, 
    8.7933, 9.4027, 7.5378, 9.2059, 19.743, 51.092, 18.875, 85.314, 62.569, 
    50.21, 82.889, 75.717, 5.5545, 0.31192, 88.296, 87.404, 16.162, 86.29, 
    4.6578, 63.086, 13.308, 23.276, 59.108, 47.609, 28.989, 74.702, 62.22, 
    26.785, 17.171, 70.991, 6.0888, 71.282, 62.54, 75.762, 60.976, 29.862, 
    37.801, 22.838, 39.681, 52.335, 7.4029, 70.28, 24.421, 93.792, 71.185, 
    77.406, 73.519, 30.726, 6.6118, 48.481, 38.466, 70.275, 41.388, 0.57959, 
    63.85, 43.84, 38.254, 93.081, 53.651, 77.428, 52.87, 13.848, 63.897, 
    89.726, 15.482, 43.941, 11.537, 73.997, 30.197, 7.8007, 60.823, 59.669, 
    27.773 ;

 alt_refrac =
  70350, 15659, 27639, 82353, 4473, 61691, 60519, 56497, 18361, 61150, 96084, 
    74349, 68875, 73030, 85964, 50499, 42939, 48674, 22200, 52846, 55785, 
    48360, 17476, 3641.6, 18145, 48263, 50894, 15042, 30638, 41919, 51411, 
    92616, 50912, 21339, 94245, 46849, 3327.8, 43829, 65451, 88280, 12151, 
    74109, 57733, 80391, 3801.4, 68964, 14225, 94028, 58186, 11954, 14500, 
    58051, 64861, 32881, 22838, 29200, 27835, 59984, 15580, 65765, 17685, 
    22038, 41886, 12348, 74348, 63985, 87119, 52305, 16393, 62091, 51899, 
    66950, 927.84, 59799, 9841.5, 46636, 93832, 5666.8, 95219, 90892, 669.32, 
    69195, 82815, 75543, -67.823, 71145, 77568, 3099.5, 50004, 97894, 82089, 
    7871.8, 77200, 46112, 74111, 10424, 45292, 10127, 37619, 55252 ;

 geop_refrac =
  8906, 22635, 37748, 2849.8, 11649, 45463, 21229, 70370, 72456, 49392, 
    40581, 25965, 90888, -103.18, 51627, 15145, 12305, 26785, 9026.2, 25975, 
    8489, 76428, 67358, 18153, 18780, 37579, 39873, 65379, 66906, 24109, 
    95822, 69880, 42301, 20917, 57095, 31686, 72587, 73898, 20038, 15407, 
    52453, 23197, 61014, 34055, 53018, 70533, 47646, 51590, 2740.8, 87979, 
    43290, 78272, 88284, 26906, 27606, 96449, 78286, 88788, 9892.1, 28179, 
    13370, 36674, 70855, 65603, 85261, 58526, 14082, 33412, 91309, 91564, 
    42519, 85976, 22869, 39777, 35197, 84936, 80970, 62288, 83336, 37315, 
    42711, 21357, 21525, 86031, 48546, 66560, 27325, 54913, 9701.8, 94115, 
    84469, 33513, 43770, 10583, 17183, 41416, 29066, 65724, 26390, 27961 ;

 refrac =
  396.75, 13.005, 124.63, 81.17, 408.53, 465.51, 326.25, 198.72, 55.582, 
    158.83, 370.99, 473.38, 183.62, 208.8, 331.85, 71.053, 133.72, 277.18, 
    156.3, 371.8, 12.207, 101.24, 388.46, 263.96, 33.888, 330.75, 378.14, 
    187.09, 60.646, 145.16, 291.01, 301.77, 82.361, 85.203, 320.83, 207.96, 
    79.092, 56.462, 344.94, 379.45, 61.239, 71.192, 410.24, 332.99, 275.14, 
    394.51, 258.2, 476.31, 470.99, 10.986, 234.78, 189.55, 464.07, 35.311, 
    384.79, 448.29, 201.29, 282.35, 211.22, 275.89, 393.46, 401.18, 411.53, 
    20.154, 139.06, 285.36, 489.65, 80.451, 294.82, 248.38, 265.3, 352.75, 
    334.94, 2.4231, 21.393, 483.19, 262.8, 265.83, 170.31, 250.9, 289.02, 
    77.282, 133.18, 481.52, 249.1, 408.17, 16.065, 442.33, 95.85, 337.2, 
    180.66, 88.151, 197.12, 167.91, 377.81, 419.47, 417.5, 45.169, 256.62, 
    115.56 ;

 refrac_sigma =
  40.938, 9.584, 32.674, 31.174, 12.197, 26.79, 48.533, 10.84, 16.077, 
    3.9628, 2.4631, 25.546, 14.843, 4.9619, 5.9381, 40.525, 13.556, 14.795, 
    9.962, 37.277, 23.435, 38.102, 0.38173, 47.913, 39.34, 38.634, 13.734, 
    16.68, 12.759, 46.149, 23.605, 9.1608, 1.322, 35.292, 46.772, 18.672, 
    20.159, 26.184, 6.4629, 27.05, 15.722, 6.6704, 40.139, 18.016, 5.9334, 
    23.303, 12.833, 33.89, 43.598, 42.983, 36.365, 11.854, 12.37, 1.8226, 
    20.737, 15.277, 35.443, 45.514, 24.109, 11.884, 45.302, 29.936, 27.032, 
    30.695, 28.406, 19.581, 46.86, 4.1301, 35.872, 20.404, 10.526, 40.916, 
    32.342, 22.988, 42.119, 26.228, 22.339, 3.4106, 33.44, 28.912, 45.12, 
    1.3641, 25.258, 29.223, 4.4311, 9.2425, 30.282, 15.152, 47.216, 23.832, 
    24.552, 16.516, 32.691, 1.548, 29.842, 33.431, 12.303, 1.1873, 25.45, 
    16.872 ;

 refrac_qual =
  33.526, 57.691, 57.57, 10.308, 41.444, 84.535, 77.027, 93.48, 9.7066, 
    63.905, 51.818, 89.765, 24.551, 97.399, 62.492, 38.389, 49.561, 10.975, 
    59.853, 55.588, 46.829, 36.46, 25.154, 10.341, 68.61, 7.2817, 10.076, 
    59.954, 62.571, 15.019, 33.389, 31.71, 80.676, 84.961, 75.278, 9.3856, 
    82.184, 41.355, 62.529, 16.014, 82.592, 87.415, 90.424, 80.337, 22.819, 
    19.264, 18.432, 26.712, 44.977, 35.402, 13.206, 25.778, 12.259, 35.851, 
    5.7019, 71.06, 16.406, 93.274, 61.747, 78.861, 2.7209, 26.029, 90.494, 
    23.634, 90.24, 4.7585, 60.05, 64.894, 25.945, 63.305, 40.654, 57.342, 
    45.944, 62.848, 22.91, 57.246, 12.911, 20.095, 64.461, 59.319, 89.253, 
    74.245, 85.363, 92.158, 57.231, 53.535, 61.349, 42.287, 86.103, 22.212, 
    38.376, 7.737, 6.3085, 36.775, 7.9917, 68.699, 43.597, 88.2, 67.973, 
    62.506 ;

 dry_temp =
  302.19, 312.76, 323.94, 160.49, 319.96, 289.74, 246.1, 311.19, 226.05, 
    154.45, 271.14, 268.13, 172.41, 293.12, 207.57, 171.41, 283.54, 335.48, 
    321.79, 231.75, 222.12, 211.39, 223.3, 207.14, 248.95, 288.7, 209.97, 
    332.04, 342.41, 303.51, 249.95, 198.49, 171.67, 187.77, 157, 174.27, 
    240.67, 244.77, 274.69, 339.79, 175.11, 280.26, 288.59, 206.15, 301.18, 
    212.64, 180.84, 171.5, 243.44, 188.77, 313.34, 281.08, 156.68, 262.28, 
    339.88, 187.76, 280.41, 309.04, 306.79, 240.56, 311.38, 282.27, 245.61, 
    281.09, 326.71, 262.56, 198.26, 165.99, 155.7, 154.55, 279.83, 223.28, 
    229.2, 206.62, 342.02, 344.44, 180.68, 265.62, 340.38, 268.41, 204.06, 
    193.04, 170.59, 274.2, 242.09, 287.77, 275.64, 183.74, 304.35, 321.28, 
    209.46, 154.61, 313.62, 179.87, 192.53, 213.45, 297.49, 187.83, 255.32, 
    307.76 ;

 dry_temp_sigma =
  32.129, 22.086, 11.61, 4.692, 37.058, 38.877, 3.6428, 46.948, 13.176, 
    23.487, 40.894, 6.1311, 7.8668, 1.1504, 27.26, 0.74814, 24.063, 13.482, 
    0.3877, 25.422, 46.669, 4.922, 12.697, 4.9421, 5.0713, 33.845, 37.191, 
    46.396, 35.048, 40.934, 13.237, 6.0026, 35.805, 43.189, 48.44, 29.257, 
    42.975, 19.31, 23.709, 39.847, 11.975, 46.622, 39.311, 3.8046, 42.305, 
    35.043, 36.229, 28.711, 0.21528, 40.391, 28.067, 34.261, 29.164, 6.3718, 
    27.78, 30.231, 34.685, 40.556, 46.155, 25.491, 31.213, 39.754, 42.886, 
    42.875, 5.5952, 24.468, 34.767, 20.404, 42.392, 0.062493, 19.581, 5.082, 
    20.013, 33.506, 0.88932, 29.119, 9.0491, 15.376, 25.492, 10.588, 8.9754, 
    33.362, 21.243, 47.485, 40.992, 25.204, 0.79696, 14.762, 38.943, 0.90196, 
    13.692, 13.018, 36.251, 27.92, 19.638, 22.563, 13.758, 31.213, 9.7472, 
    8.9637 ;

 dry_temp_qual =
  66.438, 97.241, 52.347, 15.784, 66.997, 52.739, 66.34, 56.651, 72.4, 
    60.244, 40.642, 52.152, 29.265, 42.438, 24.587, 92.709, 27.535, 0.94912, 
    34.502, 22.797, 16.247, 49.807, 23.04, 64.506, 34.525, 47.487, 52.304, 
    13.852, 48.752, 75.378, 25.293, 56.424, 80.408, 26.747, 49.826, 26.93, 
    87.247, 64.253, 16.133, 95.92, 53.585, 6.0169, 70.712, 1.7276, 66.26, 
    9.4543, 80.334, 50.551, 59.678, 48.981, 56.805, 2.8165, 44.601, 43.946, 
    92.163, 90.587, 6.1922, 21.437, 60.948, 76.072, 45.514, 38.807, 33.839, 
    87.536, 86.606, 45.766, 50.639, 34.85, 20.95, 52.68, 72.594, 79.535, 
    4.2359, 34.559, 59.729, 65.676, 27.924, 44.331, 82.55, 94.382, 47.802, 
    0.062375, 39.864, 33.202, 82.395, 41.833, 31.532, 28.673, 41.095, 44.219, 
    50.649, 84.921, 25.978, 74.037, 58.342, 72.184, 69.48, 49.69, 51.294, 
    45.464 ;

 geop =
  50220, 30959, 51163, 16211, 50268, 23460, 24649, 50710, 12326, 12271, 
    57682, 57946, 6175.7, 16899, 34064, 86795, 61194, 33597, 88651, 5037.4, 
    22774, 88124, 64865, 87040, 32370, 87510, 97269, 45370, 52411, 47115, 
    27817, 88792, 14073, 48023, 22181, 56860, 68263, 60818, 83082, 30436, 
    74202, 58694, 37125, 48201, 21202, 96356, 92845, 30954, 45499, 91001, 
    81766, 51230, 17014, 3558.4, 21493, 17489, 19698, 48505, 65072, 34925, 
    3532.9, 63443, 51021, 74143, 93282, 91521, 19106, 66941, 20969, 84179, 
    76279, 59967, 45039, 7721, 33248, 19803, 24894, 31581, 24639, 58724, 
    89672, 94397, 37262, 33630, 64830, 61745, 71027, 34331, 14157, 94102, 
    59529, 378.08, 25331, 13146, 49594, 36563, 79536, 62334, 59215, 76611 ;

 geop_sigma =
  90.86, 353.72, 372.88, 157.13, 221.19, 281.73, 298.17, 338.29, 21.264, 
    222.19, 319.19, 274.26, 255.02, 100.54, 70.989, 59.095, 329.68, 346.05, 
    264.1, 40.931, 262.03, 405.96, 451.88, 471.8, 262.86, 152.24, 67.415, 
    203.5, 101.79, 245.47, 419.15, 58.179, 431.98, 211.97, 320.34, 168.52, 
    44.535, 66.395, 454.07, 375.85, 15.491, 481.2, 419.79, 19.995, 285.03, 
    79.106, 3.7146, 360.6, 17.521, 423.82, 262.15, 112.1, 177.55, 208.44, 
    301.58, 465.78, 40.484, 297.29, 423.49, 476.82, 454.78, 233.95, 93.639, 
    239.67, 445.17, 241.77, 316, 333.54, 95.941, 113.01, 320.08, 270.42, 
    75.977, 114.25, 393.1, 98.043, 418.16, 359.81, 62.758, 53.114, 97.227, 
    258.7, 432.52, 18.565, 450.9, 339.41, 51.201, 249.43, 273.74, 370.01, 
    134.84, 34.918, 272.68, 476.11, 289.59, 302.76, 465.39, 216.08, 205.5, 
    100.79 ;

 press =
  1075.7, 47.687, 105.27, 517.94, 608.74, 513.06, 552.46, 464.55, 275.47, 
    1058.1, 218.58, 409.2, 619.18, 638.77, 773.6, 262.82, 1073.6, 1043.2, 
    168.65, 227.68, 452.03, 13.102, 16.296, 4.1717, 458.72, 188.59, 249.41, 
    623.55, 252.19, 278.43, 867.96, 1022.6, 9.661, 238.01, 783.66, 724.98, 
    324.68, 1040.7, 563.33, 985.38, 543.53, 887.25, 473.43, 886.46, 539.03, 
    382.11, 682.29, 207.4, 213.18, 1067.9, 475.73, 638.48, 792.12, 330.45, 
    569.37, 764.24, 1056.3, 633.15, 825.65, 1000.1, 442.86, 988.37, 782.72, 
    450.03, 475.24, 240.2, 725.38, 96.175, 631.49, 860.49, 527.47, 743.7, 
    106.35, 515.97, 199.41, 159.62, 664.99, 659.25, 955.8, 19.279, 162.34, 
    776.91, 981.57, 622.5, 620.56, 462.5, 21.488, 719.96, 1008.7, 614.45, 
    791.29, 154.45, 560.49, 124.44, 289.07, 298.58, 424, 573.52, 716.6, 743.15 ;

 press_sigma =
  4.3011, 4.2944, 1.9454, 3.818, 4.0523, 1.5733, 4.2951, 3.8615, 1.3226, 
    4.6903, 4.2146, 2.1357, 3.7614, 0.92314, 3.4526, 2.8509, 3.9464, 2.3158, 
    1.732, 2.2121, 3.1583, 3.1761, 1.3265, 3.3445, 3.2511, 3.5491, 0.37577, 
    3.4078, 3.9521, 0.97387, 2.774, 4.8367, 1.1509, 1.0233, 2.5405, 4.5522, 
    0.78013, 0.77319, 4.7976, 3.2789, 2.9481, 2.1322, 2.0404, 2.3067, 
    0.89876, 4.8591, 1.4481, 2.1468, 1.1597, 1.4561, 3.9742, 0.012621, 
    1.4026, 1.7998, 0.78009, 4.7506, 4.4705, 1.943, 3.0478, 0.61095, 3.3843, 
    3.9847, 1.4205, 4.616, 4.202, 4.4916, 3.3426, 1.0401, 1.346, 1.6793, 
    3.7704, 1.7594, 3.8435, 3.0079, 0.9669, 0.079072, 1.2586, 4.0481, 1.6759, 
    4.1852, 3.3387, 0.12787, 3.0876, 1.8661, 1.1005, 3.4961, 3.4066, 2.8693, 
    4.11, 2.3334, 0.78317, 3.894, 2.1639, 2.6413, 1.2497, 4.7587, 3.9345, 
    0.54979, 4.7796, 0.81147 ;

 temp =
  241.78, 168.58, 171.53, 159.21, 193.42, 325.3, 277.45, 273.82, 240.56, 
    258.41, 295.28, 172.68, 204.94, 297.09, 257.02, 186.11, 313.14, 251.48, 
    196.16, 223.02, 275.79, 276.02, 220.86, 206.94, 251.43, 160.55, 337.46, 
    254.56, 178.28, 325.18, 170.02, 150.96, 208.86, 325.24, 151.07, 297.32, 
    338.62, 334.56, 169.96, 339.95, 317.33, 170.55, 198.96, 191.98, 343.24, 
    316.21, 165.1, 266.42, 154.82, 257.12, 201.74, 312.57, 271.44, 305.09, 
    279.94, 339.19, 304.63, 327.51, 195.38, 193.4, 278.98, 331.66, 240.54, 
    308.93, 177.83, 273.85, 227.85, 186.89, 204.5, 229.08, 165.78, 164.43, 
    292.4, 289.29, 321.35, 280.35, 290.65, 314.45, 289.76, 241.6, 291.27, 
    284.69, 197.76, 324.98, 281.45, 281.92, 226.76, 324.08, 291.08, 225.72, 
    331.02, 338.7, 163.48, 214.82, 232.55, 260.94, 212.21, 241.34, 321.81, 
    282.71 ;

 temp_sigma =
  1.3651, 2.1654, 0.4244, 1.4753, 1.5546, 2.635, 2.3785, 0.67114, 3.2858, 
    2.1117, 4.1689, 4.3337, 0.43753, 1.0693, 1.3459, 0.24032, 3.7303, 0.7793, 
    4.094, 4.8291, 2.4878, 2.6886, 4.2608, 4.8708, 3.777, 3.979, 1.4373, 
    4.8237, 1.4556, 3.039, 2.0365, 1.9696, 0.067819, 1.5028, 0.012249, 2.95, 
    2.8621, 0.91488, 3.3894, 1.1224, 3.6384, 3.9009, 0.4935, 3.6333, 0.44308, 
    1.6116, 4.3707, 2.5798, 2.6742, 0.13718, 2.5596, 4.8727, 2.3961, 4.3173, 
    3.0237, 0.99647, 2.0282, 3.5077, 2.8264, 3.551, 2.0895, 4.7978, 3.0393, 
    2.9224, 0.27604, 2.3805, 1.6134, 1.0635, 4.0064, 0.06217, 2.3233, 4.3869, 
    1.2812, 2.801, 0.65008, 2.8412, 3.7793, 4.4641, 2.7033, 2.449, 3.1569, 
    4.0804, 4.3984, 0.20396, 0.68306, 1.3557, 0.7107, 1.6314, 1.9896, 
    0.06857, 2.0676, 1.9558, 1.8589, 1.8814, 1.874, 1.5042, 4.7271, 3.793, 
    3.0122, 0.87838 ;

 shum =
  21.016, 14.698, 39.667, 48.425, 47.094, 11.81, 9.5243, 28.161, 1.5937, 
    41.964, 9.7132, 47.266, 17.188, 29.861, 9.6706, 7.2319, 12.249, 30.994, 
    6.5336, 38.358, 14.12, 23.791, 1.6364, 25.788, 30.657, 18.878, 42.241, 
    28.659, 11.366, 38.238, 25.701, 14.684, 7.4148, 14.493, 23.002, 47.573, 
    25.119, 6.4788, 1.2099, 46.206, 41.205, 28.578, 45.071, 38.694, 34.961, 
    26.812, 41.417, 8.7515, 0.34124, 37.76, 47.089, 23.406, 26.403, 24.053, 
    12.305, 40.658, 46.979, 36.784, 6.1066, 8.0979, 12.075, 34.263, 19.056, 
    31.709, 26.187, 7.5544, 26.291, 39.779, 3.0894, 36.044, 12.339, 33.036, 
    16.13, 7.6296, 38.141, 6.3277, 29.245, 48.613, 18.557, 26.761, 26.589, 
    31.598, 22.926, 31.914, 9.5677, 32.861, 26.199, 18.186, 20.976, 17.492, 
    26.465, 36.557, 43.367, 31.174, 2.1797, 10.682, 32.565, 2.061, 12.723, 
    33.176 ;

 shum_sigma =
  3.4671, 0.98992, 2.6807, 3.6608, 0.33053, 0.97507, 2.2592, 1.0921, 3.8458, 
    4.2365, 4.1153, 0.073707, 3.3322, 3.1679, 3.1197, 3.1569, 4.6481, 3.2011, 
    4.6843, 1.7985, 3.0298, 0.59235, 3.2533, 4.2216, 0.58253, 1.7205, 1.7543, 
    1.5978, 4.3936, 2.1449, 3.0081, 3.6056, 4.8353, 4.1054, 1.7708, 4.6938, 
    3.3746, 4.8742, 0.221, 1.7296, 3.5965, 4.3593, 2.9675, 4.0527, 3.8452, 
    0.99896, 1.6425, 1.3386, 4.493, 1.7689, 4.2463, 3.8849, 3.9423, 3.3732, 
    2.4337, 1.6584, 2.1137, 0.92495, 3.158, 4.7958, 2.3704, 2.0595, 1.8151, 
    3.8273, 2.1804, 4.7991, 0.68643, 0.87936, 4.3972, 0.28798, 3.4645, 
    0.96895, 3.574, 3.1612, 4.5258, 3.8402, 2.687, 2.7454, 2.5255, 1.9673, 
    0.12146, 3.9996, 3.4658, 2.0884, 3.0287, 3.7486, 1.9047, 0.90397, 1.8624, 
    2.6406, 2.6956, 0.046741, 2.4122, 0.92124, 1.095, 0.67355, 3.7299, 
    0.63078, 0.052621, 0.1712 ;

 meteo_qual =
  58.231, 33.033, 82.102, 1.2224, 15.408, 87.695, 86.84, 12.26, 4.0498, 
    14.316, 92.732, 21.541, 59.203, 86.459, 18.61, 77.134, 80.209, 25.141, 
    45.814, 16.228, 95.701, 28.465, 89.794, 2.2322, 68.651, 87.156, 44.97, 
    44.973, 29.915, 92.778, 31, 69.413, 78.639, 81.767, 46.573, 73.645, 
    78.958, 17.313, 6.4881, 79.485, 9.5065, 13.939, 30.409, 74.997, 4.2438, 
    75.231, 74.437, 79.76, 61.614, 26.163, 36.935, 89.995, 55.544, 37.756, 
    49.99, 13.993, 35.795, 9.5141, 78.618, 27.19, 85.172, 93.314, 53.804, 
    41.933, 70.254, 22.451, 75.861, 82.702, 68.934, 19.204, 24.674, 69.432, 
    79.607, 53.858, 34.357, 20.614, 35.847, 28.446, 92.455, 54.556, 44.027, 
    90.415, 27.016, 69.461, 44.4, 21.902, 77.249, 18.05, 49.424, 21.391, 
    74.415, 69.788, 38.141, 62.186, 86.057, 59.736, 42.417, 77.294, 16.957, 
    47.543 ;

 geop_sfc = 5139.6 ;

 press_sfc = 669.45 ;

 press_sfc_sigma = 4.1146 ;

 press_sfc_qual = 15.749 ;

 tph_bangle = 6.2643e+06 ;

 tpa_bangle = 0.02544 ;

 tph_bangle_flag = 129 ;

 tph_refrac = 72805 ;

 tpn_refrac = 114.05 ;

 tph_refrac_flag = 56 ;

 tph_tdry_lrt = 64993 ;

 tpt_tdry_lrt = 302.82 ;

 tph_tdry_lrt_flag = 128 ;

 tph_tdry_cpt = 21745 ;

 tpt_tdry_cpt = 170.37 ;

 tph_tdry_cpt_flag = 61 ;

 prh_tdry_cpt = 28143 ;

 prt_tdry_cpt = 193.27 ;

 prh_tdry_cpt_flag = 154 ;

 tph_temp_lrt = 86692 ;

 tpt_temp_lrt = 192.36 ;

 tph_temp_lrt_flag = 107 ;

 tph_temp_cpt = 66367 ;

 tpt_temp_cpt = 316.04 ;

 tph_temp_cpt_flag = 154 ;

 prh_temp_cpt = 17682 ;

 prt_temp_cpt = 282.93 ;

 prh_temp_cpt_flag = 88 ;

 level_type =
  "METO" ;

 level_coeff_a =
  870.12, 571.26, 1306.1, 1741, 469.37, 1018.5, 629.11, 259.86, 337.9, 
    1048.6, 1820.4, 1029.5, 675.72, 703.58, 1470.6, 185.4, 840.73, 1569.9, 
    1094.9, 1785.2, 1947.1, 418.65, 313.29, 1756.3, 1628.3, 1657.5, 1346.1, 
    587.28, 375.12, 132.48, 692.47, 846.78, 1227.8, 1297.6, 1119.8, 1940.3, 
    750.49, 1376.4, 371.01, 1062.5, 249.76, 1667.6, 1624.9, 1583.2, 1617.5, 
    951.38, 1531.3, 1189.8, 419.91, 1083.6, 816.3, 88.053, 805.64, 232.34, 
    1881.8, 1480.5, 1665.7, 1672.8, 902.35, 412.06, 357.85, 747.34, 1180.6, 
    334.48, 705.17, 1148.6, 1123.1, 1218.6, 927.55, 1956.5, 1797.5, 1000.3, 
    1656.4, 488.22, 1145.4, 1578, 522.81, 1448.4, 1083.3, 868.2, 148.59, 
    749.18, 522.87, 599.83, 587.92, 1647.5, 1423.5, 42.859, 1193.2, 151.4, 
    1856.1, 403.14, 1229.3, 834.32, 781.35, 1114.5, 1185.3, 1672.3, 287.11, 
    716.4 ;

 level_coeff_b =
  1.2861, 1.102, 1.887, 1.4282, 0.42282, 0.056826, 0.1324, 0.092319, 1.2595, 
    0.11938, 1.5131, 0.99147, 1.3403, 1.4479, 1.9074, 1.4625, 0.91458, 
    1.3108, 1.0745, 0.45678, 1.6482, 1.3522, 0.52385, 0.99939, 1.5854, 
    1.3368, 0.95354, 0.8945, 0.51153, 1.7889, 0.11468, 0.028101, 1.7473, 
    0.65137, 0.68171, 0.62205, 1.3562, 1.6337, 1.8592, 0.50202, 0.035537, 
    1.1616, 0.35657, 0.0032321, 0.85188, 1.1401, 0.36367, 1.6771, 0.081564, 
    0.87803, 0.64281, 0.61784, 1.7704, 1.5729, 1.5434, 1.9251, 1.2218, 
    0.68847, 1.7756, 0.9476, 1.4298, 0.89467, 1.0152, 0.31144, 0.87682, 
    0.63174, 0.93089, 1.6374, 0.96618, 0.08647, 1.1612, 0.68791, 1.0818, 
    1.8321, 1.5034, 1.4891, 0.97672, 1.8332, 0.87081, 1.5781, 0.78089, 
    0.93451, 1.3265, 1.6935, 0.85884, 1.1886, 1.5637, 1.7367, 0.54588, 
    1.1775, 1.1907, 1.4259, 0.011319, 0.71836, 0.56175, 0.37773, 1.3616, 
    1.5212, 1.2299, 0.95752 ;
}
