netcdf ucar_testr {
dimensions:
	dim_unlim = UNLIMITED ; // (1 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1b = 5391 ;
	dim_lev2a = 5391 ;
	dim_lev2b = 5391 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 360. ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 360. ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float alt_refrac(dim_unlim, dim_lev2a) ;
		alt_refrac:long_name = "Geometric height above geoid for refractivity" ;
		alt_refrac:units = "metres" ;
		alt_refrac:valid_range = -1000., 1.e+05 ;
	float geop_refrac(dim_unlim, dim_lev2a) ;
		geop_refrac:long_name = "Geopotential height above geoid for refractivity" ;
		geop_refrac:units = "geopotential metres" ;
		geop_refrac:valid_range = -1000., 1.e+05 ;
	double refrac(dim_unlim, dim_lev2a) ;
		refrac:long_name = "Refractivity" ;
		refrac:units = "N-units" ;
		refrac:valid_range = 0., 500. ;
	double refrac_sigma(dim_unlim, dim_lev2a) ;
		refrac_sigma:long_name = "Estimated error (1-sigma) for refractivity" ;
		refrac_sigma:units = "N-units" ;
		refrac_sigma:valid_range = 0., 50. ;
	float refrac_qual(dim_unlim, dim_lev2a) ;
		refrac_qual:long_name = "Quality value for refractivity" ;
		refrac_qual:units = "percent" ;
		refrac_qual:valid_range = 0., 100. ;
	double dry_temp(dim_unlim, dim_lev2a) ;
		dry_temp:long_name = "Dry temperature" ;
		dry_temp:units = "kelvin" ;
		dry_temp:valid_range = 150., 350. ;
	double dry_temp_sigma(dim_unlim, dim_lev2a) ;
		dry_temp_sigma:long_name = "Estimated error (1-sigma) for dry temperature" ;
		dry_temp_sigma:units = "kelvin" ;
		dry_temp_sigma:valid_range = 0., 50. ;
	float dry_temp_qual(dim_unlim, dim_lev2a) ;
		dry_temp_qual:long_name = "Quality value for dry temperature" ;
		dry_temp_qual:units = "percent" ;
		dry_temp_qual:valid_range = 0., 100. ;
	float geop(dim_unlim, dim_lev2b) ;
		geop:long_name = "Geopotential height above geoid for P,T,H" ;
		geop:units = "geopotential metres" ;
		geop:valid_range = -1000., 1.e+05 ;
	float geop_sigma(dim_unlim, dim_lev2b) ;
		geop_sigma:long_name = "Estimated error (1-sigma) for geopotential height" ;
		geop_sigma:units = "geopotential metres" ;
		geop_sigma:valid_range = 0., 500. ;
	double press(dim_unlim, dim_lev2b) ;
		press:long_name = "Pressure" ;
		press:units = "hPa" ;
		press:valid_range = 0.0001, 1100. ;
	float press_sigma(dim_unlim, dim_lev2b) ;
		press_sigma:long_name = "Estimated error (1-sigma) for pressure" ;
		press_sigma:units = "hPa" ;
		press_sigma:valid_range = 0., 5. ;
	double temp(dim_unlim, dim_lev2b) ;
		temp:long_name = "Temperature" ;
		temp:units = "kelvin" ;
		temp:valid_range = 150., 350. ;
	float temp_sigma(dim_unlim, dim_lev2b) ;
		temp_sigma:long_name = "Estimated error (1-sigma) for temperature" ;
		temp_sigma:units = "kelvin" ;
		temp_sigma:valid_range = 0., 5. ;
	double shum(dim_unlim, dim_lev2b) ;
		shum:long_name = "Specific humidity" ;
		shum:units = "gram / kilogram" ;
		shum:valid_range = 0., 50. ;
	float shum_sigma(dim_unlim, dim_lev2b) ;
		shum_sigma:long_name = "Estimated  error (1-sigma) in specific humidity" ;
		shum_sigma:units = "gram / kilogram" ;
		shum_sigma:valid_range = 0., 5. ;
	float meteo_qual(dim_unlim, dim_lev2b) ;
		meteo_qual:long_name = "Quality value for meteorological data" ;
		meteo_qual:units = "percent" ;
		meteo_qual:valid_range = 0., 100. ;

// global attributes:
		:title = "ROPP Radio Occultation data" ;
		:institution = "UCAR_CDAAC" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "UCAR_CDAAC" ;
		:processing_date = "2014-11-26 10:20:26.687" ;
		:pod_method = "UNKNOWN" ;
		:phase_method = "UNKNOWN" ;
		:bangle_method = "UNKNOWN" ;
		:refrac_method = "UNKNOWN" ;
		:meteo_method = "UNKNOWN" ;
		:thin_method = "NONE (Thinning disabled) [v3.1]" ;
		:software_version = "UNKNOWN" ;
		:_FillValue = -9.9999e+07 ;
data:

 occ_id =
  "OC_20090827202208_C006_G029_UCAR" ;

 gns_id =
  "G029" ;

 leo_id =
  "C006" ;

 stn_id =
  "UNKN" ;

 start_time = 3.0472e+08 ;

 year = 2009 ;

 month = 8 ;

 day = 27 ;

 hour = 20 ;

 minute = 22 ;

 second = 8 ;

 msec = 0 ;

 pcd = 128 ;

 overall_qual = 100 ;

 time = 3.0472e+08 ;

 time_offset = 89.641 ;

 lat = -53.931 ;

 lon = -36.127 ;

 undulation = 15.31 ;

 roc = 6.3843e+06 ;

 r_coc =
  -1888.8, -4237.3, 28219 ;

 azimuth = 136.62 ;

 lat_tp =
  -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, -52.854, 
    -52.854, -52.854, -52.854, -52.855, -52.855, -52.855, -52.856, -52.856, 
    -52.856, -52.857, -52.857, -52.857, -52.858, -52.859, -52.859, -52.861, 
    -52.955, -52.955, -52.956, -52.956, -52.957, -52.957, -52.957, -52.957, 
    -52.957, -52.958, -52.958, -52.958, -53.003, -53.003, -53.003, -53.003, 
    -53.003, -53.003, -53.003, -53.003, -53.003, -53.004, -53.004, -53.004, 
    -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, 
    -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, -53.004, 
    -53.004, -53.004, -53.004, -53.005, -53.005, -53.005, -53.005, -53.005, 
    -53.005, -53.005, -53.005, -53.005, -53.005, -53.005, -53.005, -53.005, 
    -53.005, -53.005, -53.005, -53.005, -53.005, -53.006, -53.006, -53.006, 
    -53.006, -53.006, -53.006, -53.006, -53.006, -53.006, -53.006, -53.006, 
    -53.006, -53.006, -53.007, -53.007, -53.007, -53.007, -53.007, -53.007, 
    -53.007, -53.007, -53.008, -53.008, -53.008, -53.008, -53.008, -53.009, 
    -53.009, -53.042, -53.043, -53.043, -53.043, -53.044, -53.044, -53.044, 
    -53.045, -53.608, -53.609, -53.61, -53.611, -53.611, -53.612, -53.612, 
    -53.613, -53.613, -53.613, -53.614, -53.614, -53.614, -53.615, -53.615, 
    -53.615, -53.616, -53.616, -53.616, -53.616, -53.617, -53.617, -53.617, 
    -53.617, -53.618, -53.618, -53.618, -53.618, -53.618, -53.619, -53.619, 
    -53.619, -53.619, -53.619, -53.619, -53.62, -53.62, -53.62, -53.62, 
    -53.62, -53.62, -53.621, -53.621, -53.621, -53.621, -53.621, -53.621, 
    -53.621, -53.622, -53.622, -53.622, -53.622, -53.622, -53.622, -53.622, 
    -53.622, -53.623, -53.623, -53.623, -53.623, -53.623, -53.623, -53.623, 
    -53.623, -53.624, -53.624, -53.624, -53.624, -53.624, -53.624, -53.624, 
    -53.624, -53.625, -53.625, -53.625, -53.625, -53.625, -53.625, -53.625, 
    -53.625, -53.626, -53.626, -53.626, -53.626, -53.626, -53.626, -53.626, 
    -53.627, -53.627, -53.627, -53.627, -53.627, -53.627, -53.627, -53.628, 
    -53.628, -53.628, -53.628, -53.628, -53.628, -53.629, -53.629, -53.629, 
    -53.629, -53.629, -53.63, -53.63, -53.63, -53.63, -53.631, -53.631, 
    -53.631, -53.631, -53.632, -53.632, -53.632, -53.633, -53.633, -53.634, 
    -53.634, -53.635, -53.636, -53.636, -53.638, -53.64, -53.643, -53.645, 
    -53.646, -53.647, -53.649, -53.65, -53.651, -53.653, -53.654, -53.657, 
    -53.663, -53.666, -53.667, -53.669, -53.67, -53.67, -53.671, -53.672, 
    -53.673, -53.673, -53.674, -53.674, -53.675, -53.676, -53.676, -53.677, 
    -53.677, -53.678, -53.678, -53.679, -53.679, -53.679, -53.68, -53.68, 
    -53.681, -53.681, -53.682, -53.682, -53.682, -53.683, -53.683, -53.684, 
    -53.684, -53.685, -53.685, -53.685, -53.686, -53.686, -53.687, -53.71, 
    -53.712, -53.714, -53.715, -53.716, -53.717, -53.718, -53.719, -53.72, 
    -53.785, -53.785, -53.786, -53.786, -53.786, -53.786, -53.787, -53.787, 
    -53.787, -53.788, -53.788, -53.788, -53.788, -53.789, -53.789, -53.789, 
    -53.79, -53.79, -53.79, -53.791, -53.791, -53.791, -53.792, -53.792, 
    -53.792, -53.793, -53.793, -53.793, -53.794, -53.794, -53.794, -53.795, 
    -53.795, -53.795, -53.796, -53.796, -53.797, -53.797, -53.797, -53.798, 
    -53.798, -53.798, -53.799, -53.799, -53.8, -53.8, -53.8, -53.801, 
    -53.801, -53.802, -53.802, -53.802, -53.803, -53.803, -53.804, -53.804, 
    -53.805, -53.805, -53.806, -53.806, -53.807, -53.808, -53.809, -53.81, 
    -53.812, -53.817, -53.825, -53.827, -53.829, -53.83, -53.83, -53.831, 
    -53.832, -53.832, -53.833, -53.833, -53.833, -53.834, -53.834, -53.834, 
    -53.835, -53.835, -53.835, -53.836, -53.836, -53.836, -53.836, -53.837, 
    -53.837, -53.837, -53.838, -53.838, -53.838, -53.838, -53.839, -53.839, 
    -53.839, -53.839, -53.84, -53.84, -53.84, -53.84, -53.841, -53.841, 
    -53.841, -53.841, -53.842, -53.842, -53.842, -53.843, -53.843, -53.843, 
    -53.844, -53.844, -53.845, -53.845, -53.846, -53.846, -53.847, -53.847, 
    -53.848, -53.849, -53.851, -53.853, -53.855, -53.857, -53.858, -53.859, 
    -53.86, -53.861, -53.861, -53.862, -53.862, -53.863, -53.863, -53.864, 
    -53.864, -53.865, -53.865, -53.866, -53.866, -53.867, -53.867, -53.868, 
    -53.868, -53.869, -53.869, -53.87, -53.87, -53.871, -53.872, -53.959, 
    -53.96, -53.96, -53.961, -53.961, -53.961, -53.962, -53.962, -53.962, 
    -53.962, -53.962, -53.963, -53.963, -53.963, -53.963, -53.963, -53.963, 
    -53.964, -53.964, -53.964, -53.964, -53.964, -53.964, -53.964, -53.965, 
    -53.965, -53.965, -53.965, -53.965, -53.965, -53.965, -53.965, -53.966, 
    -53.966, -53.966, -53.966, -53.966, -53.966, -53.966, -53.966, -53.966, 
    -53.967, -53.967, -53.967, -53.967, -53.967, -53.967, -53.967, -53.967, 
    -53.968, -53.968, -53.968, -53.968, -53.968, -53.968, -53.968, -53.968, 
    -53.968, -53.969, -53.969, -53.969, -53.969, -53.969, -53.969, -53.969, 
    -53.969, -53.969, -53.97, -53.97, -53.97, -53.97, -53.97, -53.97, -53.97, 
    -53.97, -53.971, -53.971, -53.971, -53.971, -53.971, -53.971, -53.971, 
    -53.972, -53.972, -53.972, -53.972, -53.972, -53.972, -53.972, -53.973, 
    -53.973, -53.973, -53.973, -53.973, -53.973, -53.974, -53.974, -53.974, 
    -53.974, -53.974, -53.975, -53.975, -53.975, -53.975, -53.975, -53.975, 
    -53.976, -53.976, -53.976, -53.976, -53.976, -53.977, -53.977, -53.977, 
    -53.977, -53.977, -53.977, -53.978, -53.978, -53.978, -53.978, -53.978, 
    -53.978, -53.979, -53.979, -53.979, -53.979, -53.979, -53.979, -53.98, 
    -53.98, -53.98, -53.98, -53.98, -53.98, -53.98, -53.98, -53.981, -53.981, 
    -53.981, -53.981, -53.981, -53.981, -53.981, -53.981, -53.982, -53.982, 
    -53.982, -53.982, -53.982, -53.982, -53.982, -53.982, -53.983, -53.983, 
    -53.983, -53.983, -53.983, -53.983, -53.983, -53.983, -53.983, -53.983, 
    -53.984, -53.984, -53.984, -53.984, -53.984, -53.984, -53.984, -53.984, 
    -53.984, -53.984, -53.985, -53.985, -53.985, -53.985, -53.985, -53.985, 
    -53.985, -53.985, -53.985, -53.986, -53.986, -53.986, -53.986, -53.986, 
    -53.986, -53.986, -53.986, -53.986, -53.986, -53.987, -53.987, -53.987, 
    -53.987, -53.987, -53.987, -53.987, -53.987, -53.987, -53.987, -53.987, 
    -53.987, -53.987, -53.987, -53.988, -53.988, -53.988, -53.988, -53.988, 
    -53.988, -53.988, -53.988, -53.988, -53.988, -53.988, -53.988, -53.988, 
    -53.988, -53.988, -53.988, -53.988, -53.989, -53.989, -53.989, -53.989, 
    -53.989, -53.989, -53.989, -53.989, -53.989, -53.989, -53.989, -53.989, 
    -53.989, -53.989, -53.989, -53.99, -53.99, -53.99, -53.99, -53.99, 
    -53.99, -53.99, -53.99, -53.99, -53.99, -53.99, -53.99, -53.991, -53.991, 
    -53.991, -53.991, -53.991, -53.991, -53.991, -53.991, -53.991, -53.991, 
    -53.991, -53.991, -53.992, -53.992, -53.992, -53.992, -53.992, -53.992, 
    -53.992, -53.992, -53.992, -53.993, -53.993, -53.993, -53.993, -53.993, 
    -53.993, -53.993, -53.993, -53.994, -53.994, -53.994, -53.994, -53.994, 
    -53.994, -53.994, -53.995, -53.995, -53.995, -53.995, -53.995, -53.996, 
    -53.996, -53.996, -53.996, -53.996, -53.997, -53.997, -53.997, -53.997, 
    -53.998, -53.998, -53.998, -53.999, -53.999, -54, -54, -54.001, -54.002, 
    -54.003, -54.004, -54.006, -54.01, -54.014, -54.016, -54.018, -54.019, 
    -54.02, -54.021, -54.022, -54.023, -54.024, -54.025, -54.026, -54.027, 
    -54.028, -54.03, -54.031, -54.032, -54.033, -54.034, -54.036, -54.037, 
    -54.038, -54.039, -54.04, -54.042, -54.043, -54.044, -54.045, -54.047, 
    -54.048, -54.05, -54.053, -54.057, -54.06, -54.062, -54.063, -54.064, 
    -54.065, -54.066, -54.066, -54.067, -54.067, -54.068, -54.068, -54.069, 
    -54.069, -54.07, -54.07, -54.07, -54.071, -54.071, -54.071, -54.072, 
    -54.072, -54.072, -54.073, -54.073, -54.073, -54.074, -54.074, -54.074, 
    -54.075, -54.075, -54.075, -54.075, -54.076, -54.076, -54.076, -54.077, 
    -54.077, -54.077, -54.077, -54.078, -54.078, -54.078, -54.078, -54.079, 
    -54.079, -54.079, -54.08, -54.08, -54.08, -54.08, -54.081, -54.081, 
    -54.081, -54.082, -54.082, -54.082, -54.083, -54.083, -54.083, -54.084, 
    -54.084, -54.084, -54.085, -54.085, -54.085, -54.086, -54.086, -54.086, 
    -54.087, -54.087, -54.088, -54.088, -54.089, -54.089, -54.09, -54.09, 
    -54.091, -54.091, -54.092, -54.092, -54.093, -54.093, -54.094, -54.094, 
    -54.095, -54.095, -54.096, -54.096, -54.097, -54.097, -54.098, -54.098, 
    -54.098, -54.099, -54.099, -54.1, -54.1, -54.1, -54.101, -54.101, 
    -54.101, -54.102, -54.102, -54.102, -54.103, -54.103, -54.103, -54.104, 
    -54.104, -54.104, -54.104, -54.105, -54.105, -54.105, -54.106, -54.106, 
    -54.106, -54.106, -54.107, -54.107, -54.107, -54.107, -54.107, -54.108, 
    -54.108, -54.108, -54.108, -54.109, -54.109, -54.109, -54.109, -54.11, 
    -54.11, -54.11, -54.11, -54.11, -54.111, -54.111, -54.111, -54.111, 
    -54.112, -54.112, -54.112, -54.112, -54.112, -54.113, -54.113, -54.113, 
    -54.113, -54.113, -54.114, -54.114, -54.114, -54.114, -54.115, -54.115, 
    -54.115, -54.115, -54.116, -54.116, -54.116, -54.116, -54.117, -54.117, 
    -54.117, -54.117, -54.118, -54.118, -54.118, -54.118, -54.119, -54.119, 
    -54.119, -54.119, -54.12, -54.12, -54.12, -54.121, -54.121, -54.121, 
    -54.122, -54.122, -54.122, -54.123, -54.123, -54.124, -54.124, -54.125, 
    -54.125, -54.126, -54.126, -54.127, -54.127, -54.128, -54.128, -54.129, 
    -54.13, -54.13, -54.131, -54.131, -54.132, -54.133, -54.133, -54.134, 
    -54.134, -54.135, -54.135, -54.136, -54.136, -54.137, -54.137, -54.137, 
    -54.138, -54.138, -54.139, -54.139, -54.139, -54.14, -54.14, -54.141, 
    -54.141, -54.141, -54.142, -54.142, -54.142, -54.143, -54.143, -54.143, 
    -54.144, -54.144, -54.144, -54.144, -54.145, -54.145, -54.145, -54.146, 
    -54.146, -54.146, -54.147, -54.147, -54.147, -54.148, -54.148, -54.148, 
    -54.148, -54.149, -54.149, -54.149, -54.15, -54.15, -54.15, -54.151, 
    -54.151, -54.151, -54.152, -54.152, -54.152, -54.153, -54.153, -54.153, 
    -54.154, -54.154, -54.154, -54.155, -54.155, -54.155, -54.156, -54.156, 
    -54.156, -54.157, -54.157, -54.158, -54.158, -54.158, -54.159, -54.159, 
    -54.16, -54.16, -54.16, -54.161, -54.161, -54.162, -54.162, -54.163, 
    -54.163, -54.164, -54.164, -54.164, -54.165, -54.165, -54.166, -54.166, 
    -54.167, -54.167, -54.168, -54.168, -54.168, -54.169, -54.169, -54.17, 
    -54.17, -54.17, -54.171, -54.171, -54.172, -54.172, -54.172, -54.173, 
    -54.173, -54.173, -54.174, -54.174, -54.174, -54.175, -54.175, -54.175, 
    -54.176, -54.176, -54.176, -54.176, -54.177, -54.177, -54.177, -54.177, 
    -54.178, -54.178, -54.178, -54.179, -54.179, -54.179, -54.179, -54.18, 
    -54.18, -54.18, -54.18, -54.181, -54.181, -54.181, -54.181, -54.182, 
    -54.182, -54.182, -54.182, -54.183, -54.183, -54.183, -54.183, -54.183, 
    -54.184, -54.184, -54.184, -54.184, -54.185, -54.185, -54.185, -54.185, 
    -54.186, -54.186, -54.186, -54.186, -54.187, -54.187, -54.187, -54.187, 
    -54.187, -54.188, -54.188, -54.188, -54.188, -54.189, -54.189, -54.189, 
    -54.189, -54.19, -54.19, -54.19, -54.19, -54.191, -54.191, -54.191, 
    -54.191, -54.192, -54.192, -54.192, -54.192, -54.193, -54.193, -54.193, 
    -54.193, -54.194, -54.194, -54.194, -54.195, -54.195, -54.195, -54.195, 
    -54.196, -54.196, -54.196, -54.197, -54.197, -54.197, -54.197, -54.198, 
    -54.198, -54.198, -54.199, -54.199, -54.199, -54.2, -54.2, -54.2, 
    -54.201, -54.201, -54.201, -54.202, -54.202, -54.202, -54.203, -54.203, 
    -54.203, -54.204, -54.204, -54.204, -54.205, -54.205, -54.205, -54.206, 
    -54.206, -54.206, -54.207, -54.207, -54.207, -54.208, -54.208, -54.208, 
    -54.209, -54.209, -54.21, -54.21, -54.21, -54.211, -54.211, -54.211, 
    -54.212, -54.212, -54.212, -54.213, -54.213, -54.213, -54.214, -54.214, 
    -54.214, -54.215, -54.215, -54.215, -54.216, -54.216, -54.216, -54.217, 
    -54.217, -54.217, -54.218, -54.218, -54.218, -54.219, -54.219, -54.219, 
    -54.22, -54.22, -54.22, -54.221, -54.221, -54.221, -54.222, -54.222, 
    -54.223, -54.223, -54.223, -54.224, -54.224, -54.224, -54.225, -54.225, 
    -54.225, -54.226, -54.226, -54.227, -54.227, -54.228, -54.228, -54.228, 
    -54.229, -54.229, -54.23, -54.23, -54.231, -54.231, -54.232, -54.232, 
    -54.233, -54.233, -54.234, -54.234, -54.235, -54.235, -54.236, -54.236, 
    -54.237, -54.237, -54.238, -54.238, -54.239, -54.239, -54.24, -54.24, 
    -54.241, -54.242, -54.242, -54.243, -54.243, -54.244, -54.244, -54.245, 
    -54.245, -54.246, -54.246, -54.246, -54.247, -54.247, -54.248, -54.248, 
    -54.249, -54.249, -54.25, -54.25, -54.25, -54.251, -54.251, -54.252, 
    -54.252, -54.252, -54.253, -54.253, -54.254, -54.254, -54.254, -54.255, 
    -54.255, -54.256, -54.256, -54.256, -54.257, -54.257, -54.257, -54.258, 
    -54.258, -54.259, -54.259, -54.259, -54.26, -54.26, -54.26, -54.261, 
    -54.261, -54.261, -54.262, -54.262, -54.262, -54.263, -54.263, -54.263, 
    -54.264, -54.264, -54.264, -54.265, -54.265, -54.266, -54.266, -54.266, 
    -54.267, -54.267, -54.267, -54.268, -54.268, -54.268, -54.269, -54.269, 
    -54.269, -54.27, -54.27, -54.27, -54.271, -54.271, -54.271, -54.272, 
    -54.272, -54.272, -54.273, -54.273, -54.273, -54.274, -54.274, -54.274, 
    -54.275, -54.275, -54.275, -54.275, -54.276, -54.276, -54.276, -54.277, 
    -54.277, -54.277, -54.278, -54.278, -54.278, -54.279, -54.279, -54.279, 
    -54.279, -54.28, -54.28, -54.28, -54.281, -54.281, -54.281, -54.281, 
    -54.282, -54.282, -54.282, -54.282, -54.283, -54.283, -54.283, -54.283, 
    -54.284, -54.284, -54.284, -54.284, -54.285, -54.285, -54.285, -54.285, 
    -54.286, -54.286, -54.286, -54.286, -54.287, -54.287, -54.287, -54.287, 
    -54.288, -54.288, -54.288, -54.288, -54.288, -54.289, -54.289, -54.289, 
    -54.289, -54.29, -54.29, -54.29, -54.29, -54.291, -54.291, -54.291, 
    -54.291, -54.291, -54.292, -54.292, -54.292, -54.292, -54.293, -54.293, 
    -54.293, -54.293, -54.294, -54.294, -54.294, -54.294, -54.294, -54.295, 
    -54.295, -54.295, -54.295, -54.296, -54.296, -54.296, -54.296, -54.297, 
    -54.297, -54.297, -54.297, -54.298, -54.298, -54.298, -54.298, -54.299, 
    -54.299, -54.299, -54.299, -54.3, -54.3, -54.3, -54.3, -54.301, -54.301, 
    -54.301, -54.302, -54.302, -54.302, -54.302, -54.303, -54.303, -54.303, 
    -54.304, -54.304, -54.304, -54.304, -54.305, -54.305, -54.305, -54.306, 
    -54.306, -54.306, -54.307, -54.307, -54.307, -54.307, -54.308, -54.308, 
    -54.308, -54.309, -54.309, -54.309, -54.31, -54.31, -54.31, -54.311, 
    -54.311, -54.311, -54.312, -54.312, -54.312, -54.312, -54.313, -54.313, 
    -54.313, -54.314, -54.314, -54.314, -54.315, -54.315, -54.315, -54.316, 
    -54.316, -54.316, -54.317, -54.317, -54.317, -54.318, -54.318, -54.318, 
    -54.319, -54.319, -54.319, -54.319, -54.32, -54.32, -54.32, -54.321, 
    -54.321, -54.321, -54.322, -54.322, -54.322, -54.322, -54.323, -54.323, 
    -54.323, -54.324, -54.324, -54.324, -54.324, -54.325, -54.325, -54.325, 
    -54.325, -54.326, -54.326, -54.326, -54.327, -54.327, -54.327, -54.327, 
    -54.328, -54.328, -54.328, -54.328, -54.329, -54.329, -54.329, -54.329, 
    -54.33, -54.33, -54.33, -54.33, -54.331, -54.331, -54.331, -54.331, 
    -54.331, -54.332, -54.332, -54.332, -54.332, -54.333, -54.333, -54.333, 
    -54.333, -54.334, -54.334, -54.334, -54.334, -54.335, -54.335, -54.335, 
    -54.335, -54.336, -54.336, -54.336, -54.336, -54.337, -54.337, -54.337, 
    -54.337, -54.338, -54.338, -54.338, -54.338, -54.339, -54.339, -54.339, 
    -54.339, -54.34, -54.34, -54.34, -54.34, -54.341, -54.341, -54.341, 
    -54.342, -54.342, -54.342, -54.342, -54.343, -54.343, -54.343, -54.344, 
    -54.344, -54.344, -54.344, -54.345, -54.345, -54.345, -54.346, -54.346, 
    -54.346, -54.347, -54.347, -54.347, -54.348, -54.348, -54.348, -54.349, 
    -54.349, -54.349, -54.35, -54.35, -54.35, -54.351, -54.351, -54.351, 
    -54.352, -54.352, -54.353, -54.353, -54.353, -54.354, -54.354, -54.354, 
    -54.355, -54.355, -54.356, -54.356, -54.356, -54.357, -54.357, -54.357, 
    -54.358, -54.358, -54.359, -54.359, -54.359, -54.36, -54.36, -54.36, 
    -54.361, -54.361, -54.362, -54.362, -54.362, -54.363, -54.363, -54.363, 
    -54.364, -54.364, -54.364, -54.364, -54.365, -54.365, -54.365, -54.366, 
    -54.366, -54.366, -54.367, -54.367, -54.367, -54.367, -54.368, -54.368, 
    -54.368, -54.369, -54.369, -54.369, -54.369, -54.37, -54.37, -54.37, 
    -54.371, -54.371, -54.371, -54.371, -54.372, -54.372, -54.372, -54.372, 
    -54.373, -54.373, -54.373, -54.373, -54.374, -54.374, -54.374, -54.375, 
    -54.375, -54.375, -54.375, -54.376, -54.376, -54.376, -54.376, -54.377, 
    -54.377, -54.377, -54.377, -54.378, -54.378, -54.378, -54.379, -54.379, 
    -54.379, -54.379, -54.38, -54.38, -54.38, -54.38, -54.381, -54.381, 
    -54.381, -54.382, -54.382, -54.382, -54.382, -54.383, -54.383, -54.383, 
    -54.384, -54.384, -54.384, -54.384, -54.385, -54.385, -54.385, -54.386, 
    -54.386, -54.386, -54.386, -54.387, -54.387, -54.387, -54.388, -54.388, 
    -54.388, -54.388, -54.389, -54.389, -54.389, -54.389, -54.39, -54.39, 
    -54.39, -54.39, -54.391, -54.391, -54.391, -54.391, -54.392, -54.392, 
    -54.392, -54.392, -54.393, -54.393, -54.393, -54.393, -54.394, -54.394, 
    -54.394, -54.394, -54.395, -54.395, -54.395, -54.395, -54.396, -54.396, 
    -54.396, -54.396, -54.396, -54.397, -54.397, -54.397, -54.397, -54.397, 
    -54.398, -54.398, -54.398, -54.398, -54.398, -54.399, -54.399, -54.399, 
    -54.399, -54.399, -54.4, -54.4, -54.4, -54.4, -54.4, -54.401, -54.401, 
    -54.401, -54.401, -54.401, -54.402, -54.402, -54.402, -54.402, -54.402, 
    -54.403, -54.403, -54.403, -54.403, -54.403, -54.403, -54.404, -54.404, 
    -54.404, -54.404, -54.404, -54.405, -54.405, -54.405, -54.405, -54.405, 
    -54.406, -54.406, -54.406, -54.406, -54.406, -54.407, -54.407, -54.407, 
    -54.407, -54.407, -54.408, -54.408, -54.408, -54.408, -54.408, -54.409, 
    -54.409, -54.409, -54.409, -54.409, -54.41, -54.41, -54.41, -54.41, 
    -54.41, -54.411, -54.411, -54.411, -54.411, -54.412, -54.412, -54.412, 
    -54.412, -54.412, -54.413, -54.413, -54.413, -54.413, -54.414, -54.414, 
    -54.414, -54.415, -54.415, -54.415, -54.415, -54.416, -54.416, -54.416, 
    -54.417, -54.417, -54.417, -54.418, -54.418, -54.418, -54.419, -54.419, 
    -54.419, -54.42, -54.42, -54.42, -54.421, -54.421, -54.421, -54.422, 
    -54.422, -54.423, -54.423, -54.423, -54.424, -54.424, -54.424, -54.425, 
    -54.425, -54.426, -54.426, -54.426, -54.427, -54.427, -54.427, -54.428, 
    -54.428, -54.429, -54.429, -54.429, -54.43, -54.43, -54.43, -54.431, 
    -54.431, -54.431, -54.432, -54.432, -54.432, -54.433, -54.433, -54.433, 
    -54.433, -54.434, -54.434, -54.434, -54.435, -54.435, -54.435, -54.436, 
    -54.436, -54.436, -54.436, -54.437, -54.437, -54.437, -54.438, -54.438, 
    -54.438, -54.439, -54.439, -54.439, -54.439, -54.44, -54.44, -54.44, 
    -54.441, -54.441, -54.441, -54.441, -54.442, -54.442, -54.442, -54.443, 
    -54.443, -54.443, -54.443, -54.444, -54.444, -54.444, -54.445, -54.445, 
    -54.445, -54.446, -54.446, -54.446, -54.446, -54.447, -54.447, -54.447, 
    -54.448, -54.448, -54.448, -54.449, -54.449, -54.449, -54.449, -54.45, 
    -54.45, -54.45, -54.451, -54.451, -54.451, -54.452, -54.452, -54.452, 
    -54.453, -54.453, -54.453, -54.453, -54.454, -54.454, -54.454, -54.455, 
    -54.455, -54.455, -54.456, -54.456, -54.456, -54.456, -54.457, -54.457, 
    -54.457, -54.458, -54.458, -54.458, -54.458, -54.459, -54.459, -54.459, 
    -54.46, -54.46, -54.46, -54.46, -54.461, -54.461, -54.461, -54.462, 
    -54.462, -54.462, -54.462, -54.463, -54.463, -54.463, -54.464, -54.464, 
    -54.464, -54.464, -54.465, -54.465, -54.465, -54.465, -54.466, -54.466, 
    -54.466, -54.466, -54.467, -54.467, -54.467, -54.467, -54.468, -54.468, 
    -54.468, -54.469, -54.469, -54.469, -54.469, -54.47, -54.47, -54.47, 
    -54.47, -54.471, -54.471, -54.471, -54.471, -54.472, -54.472, -54.472, 
    -54.472, -54.473, -54.473, -54.473, -54.473, -54.474, -54.474, -54.474, 
    -54.474, -54.475, -54.475, -54.475, -54.475, -54.476, -54.476, -54.476, 
    -54.476, -54.477, -54.477, -54.477, -54.477, -54.477, -54.478, -54.478, 
    -54.478, -54.478, -54.479, -54.479, -54.479, -54.479, -54.48, -54.48, 
    -54.48, -54.48, -54.481, -54.481, -54.481, -54.481, -54.482, -54.482, 
    -54.482, -54.482, -54.483, -54.483, -54.483, -54.483, -54.484, -54.484, 
    -54.484, -54.484, -54.485, -54.485, -54.485, -54.485, -54.486, -54.486, 
    -54.486, -54.486, -54.487, -54.487, -54.487, -54.487, -54.488, -54.488, 
    -54.488, -54.488, -54.489, -54.489, -54.489, -54.489, -54.49, -54.49, 
    -54.49, -54.49, -54.491, -54.491, -54.491, -54.491, -54.492, -54.492, 
    -54.492, -54.492, -54.493, -54.493, -54.493, -54.494, -54.494, -54.494, 
    -54.494, -54.495, -54.495, -54.495, -54.495, -54.496, -54.496, -54.496, 
    -54.496, -54.497, -54.497, -54.497, -54.497, -54.498, -54.498, -54.498, 
    -54.498, -54.499, -54.499, -54.499, -54.499, -54.5, -54.5, -54.5, -54.5, 
    -54.501, -54.501, -54.501, -54.501, -54.501, -54.502, -54.502, -54.502, 
    -54.502, -54.503, -54.503, -54.503, -54.503, -54.504, -54.504, -54.504, 
    -54.504, -54.504, -54.505, -54.505, -54.505, -54.505, -54.506, -54.506, 
    -54.506, -54.506, -54.506, -54.507, -54.507, -54.507, -54.507, -54.507, 
    -54.508, -54.508, -54.508, -54.508, -54.508, -54.509, -54.509, -54.509, 
    -54.509, -54.509, -54.51, -54.51, -54.51, -54.51, -54.511, -54.511, 
    -54.511, -54.511, -54.511, -54.512, -54.512, -54.512, -54.512, -54.512, 
    -54.513, -54.513, -54.513, -54.513, -54.513, -54.514, -54.514, -54.514, 
    -54.514, -54.514, -54.514, -54.515, -54.515, -54.515, -54.515, -54.515, 
    -54.516, -54.516, -54.516, -54.516, -54.516, -54.517, -54.517, -54.517, 
    -54.517, -54.518, -54.518, -54.518, -54.518, -54.518, -54.519, -54.519, 
    -54.519, -54.519, -54.519, -54.52, -54.52, -54.52, -54.52, -54.52, 
    -54.521, -54.521, -54.521, -54.521, -54.521, -54.522, -54.522, -54.522, 
    -54.522, -54.523, -54.523, -54.523, -54.523, -54.523, -54.524, -54.524, 
    -54.524, -54.524, -54.525, -54.525, -54.525, -54.525, -54.525, -54.526, 
    -54.526, -54.526, -54.526, -54.527, -54.527, -54.527, -54.527, -54.528, 
    -54.528, -54.528, -54.528, -54.529, -54.529, -54.529, -54.529, -54.529, 
    -54.53, -54.53, -54.53, -54.531, -54.531, -54.531, -54.531, -54.532, 
    -54.532, -54.532, -54.532, -54.533, -54.533, -54.533, -54.533, -54.534, 
    -54.534, -54.534, -54.535, -54.535, -54.535, -54.535, -54.536, -54.536, 
    -54.536, -54.537, -54.537, -54.537, -54.538, -54.538, -54.538, -54.538, 
    -54.539, -54.539, -54.539, -54.54, -54.54, -54.54, -54.541, -54.541, 
    -54.541, -54.541, -54.542, -54.542, -54.542, -54.543, -54.543, -54.543, 
    -54.543, -54.544, -54.544, -54.544, -54.544, -54.545, -54.545, -54.545, 
    -54.546, -54.546, -54.546, -54.546, -54.547, -54.547, -54.547, -54.547, 
    -54.548, -54.548, -54.548, -54.548, -54.549, -54.549, -54.549, -54.549, 
    -54.549, -54.55, -54.55, -54.55, -54.55, -54.551, -54.551, -54.551, 
    -54.551, -54.551, -54.552, -54.552, -54.552, -54.552, -54.553, -54.553, 
    -54.553, -54.553, -54.553, -54.554, -54.554, -54.554, -54.554, -54.554, 
    -54.555, -54.555, -54.555, -54.555, -54.555, -54.556, -54.556, -54.556, 
    -54.556, -54.556, -54.557, -54.557, -54.557, -54.557, -54.557, -54.558, 
    -54.558, -54.558, -54.558, -54.558, -54.559, -54.559, -54.559, -54.559, 
    -54.559, -54.56, -54.56, -54.56, -54.56, -54.56, -54.561, -54.561, 
    -54.561, -54.561, -54.561, -54.562, -54.562, -54.562, -54.562, -54.562, 
    -54.563, -54.563, -54.563, -54.563, -54.563, -54.563, -54.564, -54.564, 
    -54.564, -54.564, -54.564, -54.565, -54.565, -54.565, -54.565, -54.565, 
    -54.566, -54.566, -54.566, -54.566, -54.566, -54.567, -54.567, -54.567, 
    -54.567, -54.567, -54.568, -54.568, -54.568, -54.568, -54.568, -54.568, 
    -54.569, -54.569, -54.569, -54.569, -54.569, -54.57, -54.57, -54.57, 
    -54.57, -54.57, -54.571, -54.571, -54.571, -54.571, -54.571, -54.571, 
    -54.572, -54.572, -54.572, -54.572, -54.572, -54.573, -54.573, -54.573, 
    -54.573, -54.573, -54.573, -54.574, -54.574, -54.574, -54.574, -54.574, 
    -54.575, -54.575, -54.575, -54.575, -54.575, -54.575, -54.576, -54.576, 
    -54.576, -54.576, -54.576, -54.576, -54.577, -54.577, -54.577, -54.577, 
    -54.577, -54.578, -54.578, -54.578, -54.578, -54.578, -54.578, -54.579, 
    -54.579, -54.579, -54.579, -54.579, -54.579, -54.58, -54.58, -54.58, 
    -54.58, -54.58, -54.581, -54.581, -54.581, -54.581, -54.581, -54.581, 
    -54.582, -54.582, -54.582, -54.582, -54.582, -54.583, -54.583, -54.583, 
    -54.583, -54.583, -54.583, -54.584, -54.584, -54.584, -54.584, -54.584, 
    -54.585, -54.585, -54.585, -54.585, -54.585, -54.586, -54.586, -54.586, 
    -54.586, -54.586, -54.587, -54.587, -54.587, -54.587, -54.587, -54.588, 
    -54.588, -54.588, -54.588, -54.588, -54.589, -54.589, -54.589, -54.589, 
    -54.589, -54.59, -54.59, -54.59, -54.59, -54.591, -54.591, -54.591, 
    -54.591, -54.591, -54.592, -54.592, -54.592, -54.592, -54.593, -54.593, 
    -54.593, -54.593, -54.594, -54.594, -54.594, -54.594, -54.595, -54.595, 
    -54.595, -54.595, -54.595, -54.596, -54.596, -54.596, -54.596, -54.597, 
    -54.597, -54.597, -54.597, -54.598, -54.598, -54.598, -54.598, -54.599, 
    -54.599, -54.599, -54.599, -54.6, -54.6, -54.6, -54.6, -54.601, -54.601, 
    -54.601, -54.601, -54.602, -54.602, -54.602, -54.602, -54.602, -54.603, 
    -54.603, -54.603, -54.603, -54.604, -54.604, -54.604, -54.604, -54.605, 
    -54.605, -54.605, -54.605, -54.606, -54.606, -54.606, -54.606, -54.606, 
    -54.607, -54.607, -54.607, -54.607, -54.608, -54.608, -54.608, -54.608, 
    -54.608, -54.609, -54.609, -54.609, -54.609, -54.61, -54.61, -54.61, 
    -54.61, -54.61, -54.611, -54.611, -54.611, -54.611, -54.611, -54.612, 
    -54.612, -54.612, -54.612, -54.612, -54.613, -54.613, -54.613, -54.613, 
    -54.613, -54.614, -54.614, -54.614, -54.614, -54.614, -54.614, -54.615, 
    -54.615, -54.615, -54.615, -54.615, -54.615, -54.616, -54.616, -54.616, 
    -54.616, -54.616, -54.616, -54.617, -54.617, -54.617, -54.617, -54.617, 
    -54.617, -54.618, -54.618, -54.618, -54.618, -54.618, -54.618, -54.618, 
    -54.619, -54.619, -54.619, -54.619, -54.619, -54.619, -54.619, -54.62, 
    -54.62, -54.62, -54.62, -54.62, -54.62, -54.62, -54.62, -54.621, -54.621, 
    -54.621, -54.621, -54.621, -54.621, -54.621, -54.621, -54.622, -54.622, 
    -54.622, -54.622, -54.622, -54.622, -54.622, -54.622, -54.623, -54.623, 
    -54.623, -54.623, -54.623, -54.623, -54.623, -54.623, -54.624, -54.624, 
    -54.624, -54.624, -54.624, -54.624, -54.624, -54.624, -54.624, -54.625, 
    -54.625, -54.625, -54.625, -54.625, -54.625, -54.625, -54.625, -54.625, 
    -54.626, -54.626, -54.626, -54.626, -54.626, -54.626, -54.626, -54.626, 
    -54.626, -54.627, -54.627, -54.627, -54.627, -54.627, -54.627, -54.627, 
    -54.627, -54.627, -54.628, -54.628, -54.628, -54.628, -54.628, -54.628, 
    -54.628, -54.628, -54.628, -54.628, -54.629, -54.629, -54.629, -54.629, 
    -54.629, -54.629, -54.629, -54.629, -54.629, -54.629, -54.63, -54.63, 
    -54.63, -54.63, -54.63, -54.63, -54.63, -54.63, -54.63, -54.631, -54.631, 
    -54.631, -54.631, -54.631, -54.631, -54.631, -54.631, -54.631, -54.631, 
    -54.632, -54.632, -54.632, -54.632, -54.632, -54.632, -54.632, -54.632, 
    -54.632, -54.632, -54.633, -54.633, -54.633, -54.633, -54.633, -54.633, 
    -54.633, -54.633, -54.633, -54.634, -54.634, -54.634, -54.634, -54.634, 
    -54.634, -54.634, -54.634, -54.634, -54.634, -54.635, -54.635, -54.635, 
    -54.635, -54.635, -54.635, -54.635, -54.635, -54.635, -54.636, -54.636, 
    -54.636, -54.636, -54.636, -54.636, -54.636, -54.636, -54.636, -54.636, 
    -54.637, -54.637, -54.637, -54.637, -54.637, -54.637, -54.637, -54.637, 
    -54.637, -54.638, -54.638, -54.638, -54.638, -54.638, -54.638, -54.638, 
    -54.638, -54.639, -54.639, -54.639, -54.639, -54.639, -54.639, -54.639, 
    -54.639, -54.639, -54.64, -54.64, -54.64, -54.64, -54.64, -54.64, -54.64, 
    -54.64, -54.641, -54.641, -54.641, -54.641, -54.641, -54.641, -54.641, 
    -54.641, -54.642, -54.642, -54.642, -54.642, -54.642, -54.642, -54.642, 
    -54.643, -54.643, -54.643, -54.643, -54.643, -54.643, -54.643, -54.644, 
    -54.644, -54.644, -54.644, -54.644, -54.644, -54.644, -54.645, -54.645, 
    -54.645, -54.645, -54.645, -54.645, -54.646, -54.646, -54.646, -54.646, 
    -54.646, -54.646, -54.647, -54.647, -54.647, -54.647, -54.647, -54.648, 
    -54.648, -54.648, -54.648, -54.648, -54.649, -54.649, -54.649, -54.649, 
    -54.649, -54.65, -54.65, -54.65, -54.65, -54.651, -54.651, -54.651, 
    -54.651, -54.652, -54.652, -54.652, -54.653, -54.653, -54.653, -54.653, 
    -54.654, -54.654, -54.654, -54.655, -54.655, -54.656, -54.656, -54.656, 
    -54.657, -54.657, -54.658, -54.658, -54.659, -54.659, -54.66, -54.66, 
    -54.661, -54.661, -54.662, -54.662, -54.663, -54.663, -54.664, -54.665, 
    -54.665, -54.666, -54.666, -54.667, -54.668, -54.668, -54.669, -54.669, 
    -54.67, -54.671, -54.671, -54.672, -54.673, -54.673, -54.674, -54.674, 
    -54.675, -54.676, -54.676, -54.677, -54.677, -54.678, -54.678, -54.679, 
    -54.679, -54.68, -54.68, -54.681, -54.681, -54.681, -54.682, -54.682, 
    -54.683, -54.683, -54.683, -54.684, -54.684, -54.684, -54.684, -54.685, 
    -54.685, -54.685, -54.686, -54.686, -54.686, -54.686, -54.687, -54.687, 
    -54.687, -54.687, -54.688, -54.688, -54.688, -54.688, -54.689, -54.689, 
    -54.689, -54.689, -54.69, -54.69, -54.69, -54.69, -54.69, -54.691, 
    -54.691, -54.691, -54.691, -54.692, -54.692, -54.692, -54.692, -54.692, 
    -54.693, -54.693, -54.693, -54.693, -54.693, -54.694, -54.694, -54.694, 
    -54.694, -54.694, -54.695, -54.695, -54.695, -54.695, -54.695, -54.696, 
    -54.696, -54.696, -54.696, -54.696, -54.697, -54.697, -54.697, -54.697, 
    -54.697, -54.698, -54.698, -54.698, -54.698, -54.698, -54.699, -54.699, 
    -54.699, -54.699, -54.699, -54.7, -54.7, -54.7, -54.7, -54.7, -54.7, 
    -54.701, -54.701, -54.701, -54.701, -54.701, -54.702, -54.702, -54.702, 
    -54.702, -54.702, -54.703, -54.703, -54.703, -54.703, -54.703, -54.704, 
    -54.704, -54.704, -54.704, -54.704, -54.704, -54.705, -54.705, -54.705, 
    -54.705, -54.705, -54.706, -54.706, -54.706, -54.706, -54.706, -54.706, 
    -54.707, -54.707, -54.707, -54.707, -54.707, -54.708, -54.708, -54.708, 
    -54.708, -54.708, -54.708, -54.709, -54.709, -54.709, -54.709, -54.709, 
    -54.71, -54.71, -54.71, -54.71, -54.71, -54.71, -54.711, -54.711, 
    -54.711, -54.711, -54.711, -54.711, -54.712, -54.712, -54.712, -54.712, 
    -54.712, -54.713, -54.713, -54.713, -54.713, -54.713, -54.713, -54.714, 
    -54.714, -54.714, -54.714, -54.714, -54.715, -54.715, -54.715, -54.715, 
    -54.715, -54.716, -54.716, -54.716, -54.716, -54.716, -54.717, -54.717, 
    -54.717, -54.717, -54.717, -54.718, -54.718, -54.718, -54.718, -54.718, 
    -54.719, -54.719, -54.719, -54.719, -54.719, -54.72, -54.72, -54.72, 
    -54.72, -54.721, -54.721, -54.721, -54.721, -54.722, -54.722, -54.722, 
    -54.722, -54.723, -54.723, -54.723, -54.724, -54.724, -54.724, -54.725, 
    -54.725, -54.725, -54.725, -54.726, -54.726, -54.726, -54.727, -54.727, 
    -54.727, -54.728, -54.728, -54.729, -54.729, -54.729, -54.73, -54.73, 
    -54.73, -54.731, -54.731, -54.732, -54.732, -54.732, -54.733, -54.733, 
    -54.733, -54.734, -54.734, -54.735, -54.735, -54.735, -54.736, -54.736, 
    -54.736, -54.737, -54.737, -54.737, -54.738, -54.738, -54.738, -54.739, 
    -54.739, -54.74, -54.74, -54.74, -54.741, -54.741, -54.741, -54.742, 
    -54.742, -54.742, -54.743, -54.743, -54.743, -54.744, -54.744, -54.744, 
    -54.745, -54.745, -54.745, -54.746, -54.746, -54.746, -54.747, -54.747, 
    -54.747, -54.748, -54.748, -54.748, -54.749, -54.749, -54.749, -54.75, 
    -54.75, -54.751, -54.751, -54.751, -54.752, -54.752, -54.752, -54.753, 
    -54.753, -54.754, -54.754, -54.754, -54.755, -54.755, -54.756, -54.756, 
    -54.756, -54.757, -54.757, -54.757, -54.758, -54.758, -54.759, -54.759, 
    -54.759, -54.76, -54.76, -54.761, -54.761, -54.761, -54.762, -54.762, 
    -54.762, -54.763, -54.763, -54.763, -54.764, -54.764, -54.764, -54.765, 
    -54.765, -54.765, -54.766, -54.766, -54.766, -54.767, -54.767, -54.767, 
    -54.768, -54.768, -54.768, -54.769, -54.769, -54.769, -54.77, -54.77, 
    -54.77, -54.771, -54.771, -54.771, -54.772, -54.772, -54.772, -54.773, 
    -54.773, -54.773, -54.774, -54.774, -54.774, -54.775, -54.775, -54.776, 
    -54.776, -54.776, -54.777, -54.777, -54.777, -54.778, -54.778, -54.778, 
    -54.779, -54.779, -54.779, -54.78, -54.78, -54.78, -54.781, -54.781, 
    -54.781, -54.782, -54.782, -54.782, -54.783, -54.783, -54.783, -54.784, 
    -54.784, -54.784, -54.785, -54.785, -54.785, -54.785, -54.786, -54.786, 
    -54.786, -54.787, -54.787, -54.787, -54.788, -54.788, -54.788, -54.788, 
    -54.789, -54.789, -54.789, -54.789, -54.79, -54.79, -54.79, -54.791, 
    -54.791, -54.791, -54.791, -54.792, -54.792, -54.792, -54.792, -54.793, 
    -54.793, -54.793, -54.793, -54.794, -54.794, -54.794, -54.794, -54.795, 
    -54.795, -54.795, -54.795, -54.796, -54.796, -54.796, -54.796, -54.797, 
    -54.797, -54.797, -54.797, -54.798, -54.798, -54.798, -54.798, -54.799, 
    -54.799, -54.799, -54.799, -54.8, -54.8, -54.8, -54.8, -54.801, -54.801, 
    -54.801, -54.801, -54.802, -54.802, -54.802, -54.802, -54.803, -54.803, 
    -54.803, -54.803, -54.804, -54.804, -54.804, -54.804, -54.805, -54.805, 
    -54.805, -54.805, -54.806, -54.806, -54.806, -54.806, -54.807, -54.807, 
    -54.807, -54.807, -54.808, -54.808, -54.808, -54.809, -54.809, -54.809, 
    -54.809, -54.81, -54.81, -54.81, -54.811, -54.811, -54.811, -54.812, 
    -54.812, -54.812, -54.813, -54.813, -54.813, -54.814, -54.814, -54.814, 
    -54.815, -54.815, -54.815, -54.816, -54.816, -54.817, -54.817, -54.817, 
    -54.818, -54.818, -54.818, -54.819, -54.819, -54.82, -54.82, -54.82, 
    -54.821, -54.821, -54.821, -54.822, -54.822, -54.822, -54.823, -54.823, 
    -54.823, -54.824, -54.824, -54.824, -54.825, -54.825, -54.825, -54.826, 
    -54.826, -54.826, -54.826, -54.827, -54.827, -54.827, -54.828, -54.828, 
    -54.828, -54.828, -54.829, -54.829, -54.829, -54.829, -54.83, -54.83, 
    -54.83, -54.83, -54.831, -54.831, -54.831, -54.831, -54.832, -54.832, 
    -54.832, -54.832, -54.833, -54.833, -54.833, -54.833, -54.833, -54.834, 
    -54.834, -54.834, -54.834, -54.835, -54.835, -54.835, -54.835, -54.835, 
    -54.836, -54.836, -54.836, -54.836, -54.837, -54.837, -54.837, -54.837, 
    -54.837, -54.838, -54.838, -54.838, -54.838, -54.839, -54.839, -54.839, 
    -54.839, -54.839, -54.84, -54.84, -54.84, -54.84, -54.841, -54.841, 
    -54.841, -54.841, -54.841, -54.842, -54.842, -54.842, -54.842, -54.843, 
    -54.843, -54.843, -54.844, -54.845, -54.846, -54.846, -54.847, -54.848, 
    -54.849, -54.85, -54.85, -54.851, -54.852, -54.853, -54.854, -54.855, 
    -54.855, -54.856, -54.857, -54.858, -54.859, -54.859, -54.86, -54.861, 
    -54.862, -54.863, -54.863, -54.864, -54.865, -54.866, -54.867, -54.867, 
    -54.868, -54.869, -54.87, -54.871, -54.871, -54.872, -54.873, -54.874, 
    -54.875, -54.876, -54.876, -54.877, -54.878, -54.879, -54.88, -54.88, 
    -54.881, -54.882, -54.883, -54.884, -54.884, -54.885, -54.886, -54.887, 
    -54.888, -54.888, -54.889, -54.89, -54.891, -54.892, -54.892, -54.893, 
    -54.894, -54.895, -54.896, -54.897, -54.897, -54.898, -54.899, -54.9, 
    -54.901, -54.901, -54.902, -54.903, -54.904, -54.905, -54.905, -54.906, 
    -54.907, -54.908, -54.909, -54.909, -54.91, -54.911, -54.912, -54.913, 
    -54.913, -54.914, -54.915, -54.916, -54.917, -54.917, -54.918, -54.919, 
    -54.92, -54.921, -54.921, -54.922, -54.923, -54.924, -54.925, -54.925, 
    -54.926, -54.927, -54.928, -54.929, -54.929, -54.93, -54.931, -54.932, 
    -54.933, -54.933, -54.934, -54.935, -54.936, -54.937, -54.937, -54.938, 
    -54.939, -54.94, -54.941, -54.941, -54.942, -54.943, -54.944, -54.945, 
    -54.945, -54.946, -54.947, -54.948, -54.949, -54.949, -54.95, -54.951, 
    -54.952, -54.953, -54.953, -54.954, -54.955, -54.956, -54.957, -54.957, 
    -54.958, -54.959, -54.96, -54.961, -54.961, -54.962, -54.963, -54.964, 
    -54.965, -54.965, -54.966, -54.967, -54.968, -54.969, -54.969, -54.97, 
    -54.971, -54.972, -54.972, -54.973, -54.974, -54.975, -54.976, -54.976, 
    -54.977, -54.978, -54.979, -54.98, -54.98, -54.981, -54.982, -54.983, 
    -54.983, -54.984, -54.985, -54.986, -54.987, -54.987, -54.988, -54.989, 
    -54.99, -54.991, -54.991, -54.992, -54.993, -54.994, -54.994, -54.995, 
    -54.996, -54.997, -54.998, -54.998, -54.999, -55, -55.001, -55.002, 
    -55.002, -55.003, -55.004, -55.005, -55.005, -55.006, -55.007, -55.008, 
    -55.009, -55.009, -55.01, -55.011, -55.012, -55.012, -55.013, -55.014, 
    -55.015, -55.016, -55.016, -55.017, -55.018, -55.019, -55.019, -55.02, 
    -55.021, -55.022, -55.022, -55.023, -55.024, -55.025, -55.025, -55.026, 
    -55.027, -55.028, -55.028, -55.029, -55.03, -55.031, -55.032, -55.032, 
    -55.033, -55.034, -55.035, -55.035, -55.036, -55.037, -55.038, -55.038, 
    -55.039, -55.04, -55.041, -55.041, -55.042, -55.043, -55.044, -55.044, 
    -55.045, -55.046, -55.047, -55.048, -55.048, -55.049, -55.05, -55.051, 
    -55.051, -55.052, -55.053, -55.054, -55.055, -55.055, -55.056, -55.057, 
    -55.058, -55.058, -55.059, -55.06, -55.061, -55.062, -55.062, -55.063, 
    -55.064, -55.065, -55.066, -55.066, -55.067, -55.068, -55.069, -55.069, 
    -55.07, -55.071, -55.072, -55.073, -55.073, -55.074, -55.075, -55.076, 
    -55.077, -55.077, -55.078, -55.079, -55.08, -55.08, -55.081, -55.082, 
    -55.083, -55.084, -55.084, -55.085, -55.086, -55.087, -55.087, -55.088, 
    -55.089, -55.09, -55.091, -55.091, -55.092, -55.093, -55.094, -55.094, 
    -55.095, -55.096, -55.097, -55.097, -55.098, -55.099, -55.1, -55.1, 
    -55.101, -55.102, -55.103, -55.103, -55.104, -55.105, -55.106, -55.106, 
    -55.107, -55.108, -55.109, -55.109, -55.11, -55.111, -55.112, -55.112, 
    -55.113, -55.114, -55.115, -55.115, -55.116, -55.117, -55.118, -55.118, 
    -55.119, -55.12, -55.121, -55.121, -55.122, -55.123, -55.124, -55.124, 
    -55.125, -55.126, -55.127, -55.127, -55.128, -55.129, -55.13, -55.13, 
    -55.131, -55.132, -55.133, -55.133, -55.134, -55.135, -55.136, -55.136, 
    -55.137, -55.138, -55.139, -55.14, -55.14, -55.141, -55.142, -55.143, 
    -55.143, -55.144, -55.145, -55.146, -55.146, -55.147, -55.148, -55.149, 
    -55.149, -55.15, -55.151, -55.152, -55.153, -55.153, -55.154, -55.155, 
    -55.156, -55.156, -55.157, -55.158, -55.159, -55.159, -55.16, -55.161, 
    -55.162, -55.162, -55.163, -55.164, -55.165, -55.165, -55.166, -55.167, 
    -55.168, -55.168, -55.169, -55.17, -55.171, -55.171, -55.172, -55.173, 
    -55.174, -55.174, -55.175, -55.176, -55.177, -55.177, -55.178, -55.179, 
    -55.18, -55.18, -55.181, -55.182, -55.183, -55.183, -55.184, -55.185, 
    -55.186, -55.186, -55.187, -55.188, -55.189, -55.189, -55.19, -55.191, 
    -55.192, -55.192, -55.193, -55.194, -55.195, -55.195, -55.196, -55.197, 
    -55.198, -55.198, -55.199, -55.2, -55.201, -55.201, -55.202, -55.203, 
    -55.204, -55.204, -55.205, -55.206, -55.207, -55.207, -55.208, -55.209, 
    -55.209, -55.21, -55.211, -55.212, -55.212, -55.213, -55.214, -55.215, 
    -55.215, -55.216, -55.217, -55.217, -55.218, -55.219, -55.22, -55.22, 
    -55.221, -55.222, -55.222, -55.223, -55.224, -55.225, -55.225, -55.226, 
    -55.227, -55.228, -55.228, -55.229, -55.23, -55.231, -55.231, -55.232, 
    -55.233, -55.234, -55.234, -55.235, -55.236, -55.236, -55.237, -55.238, 
    -55.239, -55.239, -55.24, -55.241, -55.242, -55.242, -55.243, -55.244, 
    -55.245, -55.245, -55.246, -55.247, -55.248, -55.248, -55.249, -55.25, 
    -55.251, -55.251, -55.252, -55.253, -55.253, -55.254, -55.255, -55.256, 
    -55.256, -55.257, -55.258, -55.258, -55.259, -55.26, -55.261, -55.261, 
    -55.262, -55.263, -55.263, -55.264, -55.265, -55.266, -55.266, -55.267, 
    -55.268, -55.268, -55.269, -55.27, -55.271, -55.271, -55.272, -55.273, 
    -55.273, -55.274, -55.275, -55.276, -55.276, -55.277, -55.278, -55.278, 
    -55.279, -55.28, -55.281, -55.281, -55.282, -55.283, -55.284, -55.284, 
    -55.285, -55.286, -55.286, -55.287, -55.288, -55.289, -55.289, -55.29, 
    -55.291, -55.292, -55.292, -55.293, -55.294, -55.294, -55.295, -55.296, 
    -55.297, -55.297, -55.298, -55.299, -55.3, -55.3, -55.301, -55.302, 
    -55.302, -55.303, -55.304, -55.305, -55.305, -55.306, -55.307, -55.307, 
    -55.308, -55.309, -55.309, -55.31, -55.311, -55.312, -55.312, -55.313, 
    -55.314, -55.314, -55.315, -55.316, -55.316, -55.317, -55.318, -55.319, 
    -55.319, -55.32, -55.321, -55.321, -55.322, -55.323, -55.323, -55.324, 
    -55.325, -55.326, -55.326, -55.327, -55.328, -55.328, -55.329, -55.33, 
    -55.33, -55.331, -55.332, -55.333, -55.333, -55.334, -55.335, -55.335, 
    -55.336, -55.337, -55.337, -55.338, -55.339, -55.34, -55.34, -55.341, 
    -55.342, -55.342, -55.343, -55.344, -55.345, -55.345, -55.346, -55.347, 
    -55.347, -55.348, -55.349, -55.349, -55.35, -55.351, -55.352, -55.352, 
    -55.353, -55.354, -55.354, -55.355, -55.356, -55.357, -55.357, -55.358, 
    -55.359, -55.359, -55.36, -55.361, -55.361, -55.362, -55.363, -55.364, 
    -55.364, -55.365, -55.366, -55.366, -55.367, -55.368, -55.368, -55.369, 
    -55.37, -55.371, -55.371, -55.372, -55.373, -55.373, -55.374, -55.375, 
    -55.375, -55.376, -55.377, -55.377, -55.378, -55.379, -55.379, -55.38, 
    -55.381, -55.381, -55.382, -55.383, -55.383, -55.384, -55.385, -55.386, 
    -55.386, -55.387, -55.388, -55.388, -55.389, -55.39, -55.39, -55.391, 
    -55.392, -55.392, -55.393, -55.394, -55.394, -55.395, -55.396, -55.397, 
    -55.397, -55.398, -55.399, -55.399, -55.4, -55.401, -55.401, -55.402, 
    -55.403, -55.403, -55.404, -55.405, -55.405, -55.406, -55.407, -55.408, 
    -55.408, -55.409, -55.41, -55.41, -55.411, -55.412, -55.412, -55.413, 
    -55.414, -55.414, -55.415, -55.416, -55.416, -55.417, -55.418, -55.419, 
    -55.419, -55.42, -55.421, -55.421, -55.422, -55.423, -55.423, -55.424, 
    -55.425, -55.425, -55.426, -55.427, -55.427, -55.428, -55.429, -55.43, 
    -55.43, -55.431, -55.432, -55.432, -55.433, -55.434, -55.434, -55.435, 
    -55.436, -55.436, -55.437, -55.438, -55.438, -55.439, -55.44, -55.441, 
    -55.441, -55.442, -55.443, -55.443, -55.444, -55.445, -55.445, -55.446, 
    -55.447, -55.447, -55.448, -55.449, -55.449, -55.45, -55.451, -55.451, 
    -55.452, -55.453, -55.453, -55.454, -55.455, -55.455, -55.456, -55.457, 
    -55.457, -55.458, -55.459, -55.459, -55.46, -55.461, -55.461, -55.462, 
    -55.463, -55.463, -55.464, -55.465, -55.465, -55.466, -55.467, -55.467, 
    -55.468, -55.469, -55.469, -55.47, -55.471, -55.472, -55.472, -55.473, 
    -55.474, -55.474, -55.475, -55.476, -55.476, -55.477, -55.478, -55.478, 
    -55.479, -55.48, -55.48, -55.481, -55.482, -55.482, -55.483, -55.484, 
    -55.484, -55.485, -55.486, -55.486, -55.487, -55.488, -55.488, -55.489, 
    -55.49, -55.49, -55.491, -55.492, -55.492, -55.493, -55.494, -55.494, 
    -55.495, -55.496, -55.496, -55.497, -55.498, -55.498, -55.499, -55.5, 
    -55.5, -55.501, -55.502, -55.502, -55.503, -55.504, -55.504, -55.505, 
    -55.506, -55.506, -55.507, -55.508, -55.508, -55.509, -55.51, -55.51, 
    -55.511, -55.512, -55.512, -55.513, -55.514, -55.514, -55.515, -55.516, 
    -55.516, -55.517, -55.518, -55.518, -55.519, -55.52, -55.52, -55.521, 
    -55.522, -55.522, -55.523, -55.524, -55.524, -55.525, -55.526, -55.526, 
    -55.527, -55.528, -55.528, -55.529, -55.53, -55.53, -55.531, -55.532, 
    -55.532, -55.533, -55.534, -55.534, -55.535, -55.536, -55.536, -55.537, 
    -55.538, -55.538, -55.539, -55.54, -55.54, -55.541, -55.542, -55.542, 
    -55.543, -55.544, -55.544, -55.545, -55.546, -55.546, -55.547, -55.548, 
    -55.548, -55.549, -55.55, -55.55, -55.551, -55.552, -55.552, -55.553, 
    -55.554, -55.554, -55.555, -55.556, -55.556, -55.557, -55.558, -55.558, 
    -55.559, -55.559, -55.56, -55.561, -55.561, -55.562, -55.563, -55.563, 
    -55.564, -55.565, -55.565, -55.566, -55.567, -55.567, -55.568, -55.569, 
    -55.569, -55.57, -55.571, -55.571, -55.572, -55.573, -55.573, -55.574, 
    -55.575, -55.575, -55.576, -55.577, -55.577, -55.578, -55.579, -55.579, 
    -55.58, -55.581, -55.581, -55.582, -55.583, -55.583, -55.584, -55.585, 
    -55.585, -55.586, -55.587, -55.587, -55.588, -55.589, -55.589, -55.59, 
    -55.591, -55.591, -55.592, -55.593, -55.593, -55.594, -55.595, -55.595, 
    -55.596, -55.597, -55.597, -55.598, -55.599, -55.599, -55.6, -55.601, 
    -55.601, -55.602, -55.602, -55.603, -55.604, -55.604, -55.605, -55.606, 
    -55.606, -55.607, -55.608, -55.608, -55.609, -55.61, -55.61, -55.611, 
    -55.612, -55.612, -55.613, -55.614, -55.614, -55.615, -55.616, -55.616, 
    -55.617, -55.618, -55.618, -55.619, -55.62, -55.62, -55.621, -55.622, 
    -55.622, -55.623, -55.624, -55.624, -55.625, -55.626, -55.626, -55.627, 
    -55.628, -55.628, -55.629, -55.63, -55.63, -55.631, -55.631, -55.632, 
    -55.633, -55.633, -55.634, -55.635, -55.635, -55.636, -55.637, -55.637, 
    -55.638, -55.639, -55.639, -55.64, -55.641, -55.641, -55.642, -55.643, 
    -55.643, -55.644, -55.645, -55.645, -55.646, -55.647, -55.647, -55.648, 
    -55.649, -55.649, -55.65, -55.651, -55.651, -55.652, -55.653, -55.653, 
    -55.654, -55.655, -55.655, -55.656, -55.656, -55.657, -55.658, -55.658, 
    -55.659, -55.66, -55.66, -55.661, -55.662, -55.662, -55.663, -55.664, 
    -55.664, -55.665, -55.666, -55.666, -55.667, -55.668, -55.668, -55.669, 
    -55.67, -55.67, -55.671, -55.672, -55.672, -55.673, -55.674, -55.674, 
    -55.675, -55.676, -55.676, -55.677, -55.677, -55.678, -55.679, -55.679, 
    -55.68, -55.681, -55.681, -55.682, -55.683, -55.683, -55.684, -55.685, 
    -55.685, -55.686, -55.687, -55.687, -55.688, -55.689, -55.689, -55.69, 
    -55.691, -55.691, -55.692, -55.693, -55.693, -55.694, -55.694, -55.695, 
    -55.696, -55.696, -55.697, -55.698, -55.698, -55.699, -55.7, -55.7, 
    -55.701, -55.702, -55.702, -55.703, -55.704, -55.704, -55.705, -55.706, 
    -55.706, -55.707, -55.708, -55.708, -55.709, -55.71, -55.71, -55.711, 
    -55.711, -55.712, -55.713, -55.713, -55.714, -55.715, -55.715, -55.716, 
    -55.717, -55.717, -55.718, -55.719, -55.719, -55.72, -55.721, -55.721, 
    -55.722, -55.723, -55.723, -55.724, -55.725, -55.725, -55.726, -55.727, 
    -55.727, -55.728, -55.729, -55.729, -55.73, -55.731, -55.731, -55.732, 
    -55.733, -55.733, -55.734, -55.734, -55.735, -55.736, -55.736, -55.737, 
    -55.738, -55.738, -55.739, -55.74, -55.74, -55.741, -55.742, -55.742, 
    -55.743, -55.744, -55.744, -55.745, -55.746, -55.746, -55.747, -55.747, 
    -55.748, -55.749, -55.749, -55.75, -55.751, -55.751, -55.752, -55.753, 
    -55.753, -55.754, -55.755, -55.755, -55.756, -55.757, -55.757, -55.758, 
    -55.759, -55.759, -55.76, -55.761, -55.761, -55.762, -55.763, -55.763, 
    -55.764, -55.765, -55.765, -55.766, -55.767, -55.767, -55.768, -55.768, 
    -55.769, -55.77, -55.77, -55.771, -55.772, -55.772, -55.773, -55.774, 
    -55.774, -55.775, -55.776, -55.776, -55.777, -55.778, -55.778, -55.779, 
    -55.78, -55.78, -55.781, -55.782, -55.782, -55.783, -55.784, -55.784, 
    -55.785, -55.786, -55.786, -55.787, -55.787, -55.788, -55.789, -55.789, 
    -55.79, -55.791, -55.791, -55.792, -55.793, -55.793, -55.794, -55.795, 
    -55.795, -55.796, -55.797, -55.797, -55.798, -55.799, -55.799, -55.8, 
    -55.8, -55.801, -55.802, -55.802, -55.803, -55.804, -55.804, -55.805, 
    -55.806, -55.806, -55.807, -55.808, -55.808, -55.809, -55.81, -55.81, 
    -55.811, -55.812, -55.812, -55.813, -55.814, -55.814, -55.815, -55.815, 
    -55.816, -55.817, -55.817, -55.818, -55.819, -55.819, -55.82, -55.821, 
    -55.821, -55.822, -55.823, -55.823, -55.824, -55.825, -55.825, -55.826, 
    -55.827, -55.827, -55.828, -55.829, -55.829, -55.83, -55.831, -55.831, 
    -55.832, -55.833, -55.833, -55.834, -55.835, -55.835, -55.836, -55.836, 
    -55.837, -55.838, -55.838, -55.839, -55.84, -55.84, -55.841, -55.842, 
    -55.842, -55.843, -55.844, -55.844, -55.845, -55.846, -55.846, -55.847, 
    -55.848, -55.848, -55.849, -55.85, -55.85, -55.851, -55.852, -55.852, 
    -55.853, -55.854, -55.854, -55.855, -55.856, -55.856, -55.857, -55.858, 
    -55.858, -55.859, -55.859, -55.86, -55.861, -55.861, -55.862, -55.863, 
    -55.863, -55.864, -55.865, -55.865, -55.866, -55.867, -55.867, -55.868, 
    -55.869, -55.869, -55.87, -55.871, -55.871, -55.872, -55.873, -55.873, 
    -55.874, -55.874, -55.875, -55.876, -55.876, -55.877, -55.878, -55.878, 
    -55.879, -55.88, -55.88, -55.881, -55.882, -55.882, -55.883, -55.884, 
    -55.884, -55.885, -55.886, -55.886, -55.887, -55.888, -55.888, -55.889, 
    -55.89, -55.89, -55.891, -55.891, -55.892, -55.893, -55.893, -55.894, 
    -55.895, -55.895, -55.896, -55.897, -55.897, -55.898, -55.899, -55.899, 
    -55.9, -55.901, -55.901, -55.902, -55.903, -55.903, -55.904, -55.905, 
    -55.905, -55.906, -55.907, -55.907, -55.908, -55.908, -55.909, -55.91, 
    -55.91, -55.911, -55.912, -55.912, -55.913, -55.914, -55.914, -55.915, 
    -55.916, -55.916, -55.917, -55.918, -55.918, -55.919, -55.92, -55.92, 
    -55.921, -55.922, -55.922, -55.923, -55.923, -55.924, -55.925, -55.925, 
    -55.926, -55.927, -55.927, -55.928, -55.929, -55.929, -55.93, -55.931, 
    -55.931, -55.932, -55.933, -55.933, -55.934, -55.935, -55.935, -55.936, 
    -55.936, -55.937, -55.938, -55.938, -55.939, -55.94, -55.94, -55.941, 
    -55.942, -55.942, -55.943, -55.944, -55.944, -55.945, -55.946, -55.946, 
    -55.947, -55.948, -55.948, -55.949, -55.95, -55.95, -55.951, -55.952, 
    -55.952, -55.953, -55.954, -55.954, -55.955, -55.955, -55.956, -55.957, 
    -55.957, -55.958, -55.959, -55.959, -55.96, -55.961, -55.961, -55.962, 
    -55.963, -55.963, -55.964, -55.965, -55.965, -55.966, -55.967, -55.967, 
    -55.968, -55.969, -55.969, -55.97, -55.97, -55.971, -55.972, -55.972, 
    -55.973, -55.974 ;

 lon_tp =
  -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, -35.566, 
    -35.566, -35.566, -35.566, -35.566, -35.566, -35.567, -35.567, -35.567, 
    -35.567, -35.568, -35.568, -35.568, -35.569, -35.569, -35.569, -35.57, 
    -35.606, -35.607, -35.607, -35.607, -35.608, -35.608, -35.608, -35.608, 
    -35.608, -35.609, -35.609, -35.609, -35.643, -35.643, -35.643, -35.643, 
    -35.643, -35.643, -35.644, -35.644, -35.644, -35.644, -35.644, -35.644, 
    -35.644, -35.644, -35.644, -35.644, -35.644, -35.645, -35.645, -35.645, 
    -35.645, -35.645, -35.645, -35.645, -35.645, -35.645, -35.645, -35.646, 
    -35.646, -35.646, -35.646, -35.646, -35.646, -35.646, -35.646, -35.646, 
    -35.646, -35.646, -35.647, -35.647, -35.647, -35.647, -35.647, -35.647, 
    -35.647, -35.647, -35.647, -35.647, -35.648, -35.648, -35.648, -35.648, 
    -35.648, -35.648, -35.648, -35.648, -35.648, -35.649, -35.649, -35.649, 
    -35.649, -35.649, -35.649, -35.649, -35.649, -35.649, -35.65, -35.65, 
    -35.65, -35.65, -35.65, -35.65, -35.65, -35.651, -35.651, -35.651, 
    -35.651, -35.652, -35.652, -35.652, -35.653, -35.653, -35.653, -35.653, 
    -35.654, -35.943, -35.944, -35.944, -35.945, -35.945, -35.945, -35.946, 
    -35.946, -35.946, -35.947, -35.947, -35.947, -35.947, -35.948, -35.948, 
    -35.948, -35.948, -35.949, -35.949, -35.949, -35.949, -35.949, -35.95, 
    -35.95, -35.95, -35.95, -35.95, -35.95, -35.951, -35.951, -35.951, 
    -35.951, -35.951, -35.951, -35.952, -35.952, -35.952, -35.952, -35.952, 
    -35.952, -35.953, -35.953, -35.953, -35.953, -35.953, -35.953, -35.953, 
    -35.954, -35.954, -35.954, -35.954, -35.954, -35.954, -35.954, -35.954, 
    -35.955, -35.955, -35.955, -35.955, -35.955, -35.955, -35.955, -35.956, 
    -35.956, -35.956, -35.956, -35.956, -35.956, -35.956, -35.957, -35.957, 
    -35.957, -35.957, -35.957, -35.957, -35.957, -35.957, -35.958, -35.958, 
    -35.958, -35.958, -35.958, -35.958, -35.958, -35.959, -35.959, -35.959, 
    -35.959, -35.959, -35.959, -35.959, -35.96, -35.96, -35.96, -35.96, 
    -35.96, -35.96, -35.961, -35.961, -35.961, -35.961, -35.961, -35.961, 
    -35.961, -35.962, -35.962, -35.962, -35.962, -35.962, -35.963, -35.963, 
    -35.963, -35.963, -35.963, -35.964, -35.964, -35.964, -35.965, -35.965, 
    -35.965, -35.966, -35.966, -35.967, -35.967, -35.969, -35.97, -35.971, 
    -35.972, -35.973, -35.973, -35.974, -35.975, -35.976, -35.977, -35.978, 
    -35.981, -35.983, -35.984, -35.984, -35.985, -35.985, -35.986, -35.986, 
    -35.987, -35.987, -35.988, -35.988, -35.988, -35.989, -35.989, -35.989, 
    -35.99, -35.99, -35.99, -35.991, -35.991, -35.991, -35.992, -35.992, 
    -35.992, -35.992, -35.993, -35.993, -35.993, -35.994, -35.994, -35.994, 
    -35.994, -35.995, -35.995, -35.995, -35.996, -35.996, -35.997, -36.008, 
    -36.009, -36.01, -36.011, -36.012, -36.012, -36.013, -36.013, -36.014, 
    -36.051, -36.051, -36.051, -36.052, -36.052, -36.052, -36.052, -36.052, 
    -36.053, -36.053, -36.053, -36.053, -36.054, -36.054, -36.054, -36.054, 
    -36.054, -36.055, -36.055, -36.055, -36.055, -36.056, -36.056, -36.056, 
    -36.056, -36.057, -36.057, -36.057, -36.057, -36.058, -36.058, -36.058, 
    -36.058, -36.059, -36.059, -36.059, -36.059, -36.06, -36.06, -36.06, 
    -36.061, -36.061, -36.061, -36.061, -36.062, -36.062, -36.062, -36.062, 
    -36.063, -36.063, -36.063, -36.064, -36.064, -36.064, -36.064, -36.065, 
    -36.065, -36.065, -36.066, -36.066, -36.067, -36.067, -36.068, -36.069, 
    -36.07, -36.072, -36.076, -36.078, -36.078, -36.079, -36.079, -36.08, 
    -36.08, -36.081, -36.081, -36.081, -36.081, -36.082, -36.082, -36.082, 
    -36.082, -36.083, -36.083, -36.083, -36.083, -36.084, -36.084, -36.084, 
    -36.084, -36.084, -36.085, -36.085, -36.085, -36.085, -36.085, -36.086, 
    -36.086, -36.086, -36.086, -36.086, -36.087, -36.087, -36.087, -36.087, 
    -36.087, -36.088, -36.088, -36.088, -36.088, -36.089, -36.089, -36.089, 
    -36.089, -36.09, -36.09, -36.09, -36.091, -36.091, -36.091, -36.092, 
    -36.092, -36.093, -36.094, -36.095, -36.096, -36.097, -36.098, -36.098, 
    -36.099, -36.099, -36.1, -36.1, -36.1, -36.101, -36.101, -36.102, 
    -36.102, -36.102, -36.102, -36.103, -36.103, -36.103, -36.104, -36.104, 
    -36.104, -36.105, -36.105, -36.105, -36.106, -36.106, -36.107, -36.138, 
    -36.139, -36.139, -36.139, -36.139, -36.14, -36.14, -36.14, -36.14, 
    -36.14, -36.141, -36.141, -36.141, -36.141, -36.141, -36.141, -36.142, 
    -36.142, -36.142, -36.142, -36.142, -36.142, -36.142, -36.143, -36.143, 
    -36.143, -36.143, -36.143, -36.143, -36.143, -36.144, -36.144, -36.144, 
    -36.144, -36.144, -36.144, -36.144, -36.144, -36.145, -36.145, -36.145, 
    -36.145, -36.145, -36.145, -36.145, -36.146, -36.146, -36.146, -36.146, 
    -36.146, -36.146, -36.146, -36.146, -36.147, -36.147, -36.147, -36.147, 
    -36.147, -36.147, -36.147, -36.147, -36.148, -36.148, -36.148, -36.148, 
    -36.148, -36.148, -36.148, -36.149, -36.149, -36.149, -36.149, -36.149, 
    -36.149, -36.149, -36.149, -36.15, -36.15, -36.15, -36.15, -36.15, 
    -36.15, -36.15, -36.151, -36.151, -36.151, -36.151, -36.151, -36.151, 
    -36.152, -36.152, -36.152, -36.152, -36.152, -36.152, -36.153, -36.153, 
    -36.153, -36.153, -36.153, -36.153, -36.153, -36.154, -36.154, -36.154, 
    -36.154, -36.154, -36.154, -36.155, -36.155, -36.155, -36.155, -36.155, 
    -36.155, -36.156, -36.156, -36.156, -36.156, -36.156, -36.156, -36.157, 
    -36.157, -36.157, -36.157, -36.157, -36.157, -36.158, -36.158, -36.158, 
    -36.158, -36.158, -36.158, -36.158, -36.159, -36.159, -36.159, -36.159, 
    -36.159, -36.159, -36.159, -36.16, -36.16, -36.16, -36.16, -36.16, 
    -36.16, -36.16, -36.16, -36.161, -36.161, -36.161, -36.161, -36.161, 
    -36.161, -36.161, -36.161, -36.162, -36.162, -36.162, -36.162, -36.162, 
    -36.162, -36.162, -36.163, -36.163, -36.163, -36.163, -36.163, -36.163, 
    -36.163, -36.163, -36.164, -36.164, -36.164, -36.164, -36.164, -36.164, 
    -36.164, -36.164, -36.164, -36.165, -36.165, -36.165, -36.165, -36.165, 
    -36.165, -36.165, -36.165, -36.166, -36.166, -36.166, -36.166, -36.166, 
    -36.166, -36.166, -36.166, -36.167, -36.167, -36.167, -36.167, -36.167, 
    -36.167, -36.167, -36.167, -36.167, -36.167, -36.167, -36.167, -36.167, 
    -36.167, -36.167, -36.168, -36.168, -36.168, -36.168, -36.168, -36.168, 
    -36.168, -36.168, -36.168, -36.168, -36.168, -36.168, -36.168, -36.168, 
    -36.169, -36.169, -36.169, -36.169, -36.169, -36.169, -36.169, -36.169, 
    -36.169, -36.169, -36.169, -36.169, -36.169, -36.169, -36.17, -36.17, 
    -36.17, -36.17, -36.17, -36.17, -36.17, -36.17, -36.17, -36.17, -36.17, 
    -36.17, -36.17, -36.171, -36.171, -36.171, -36.171, -36.171, -36.171, 
    -36.171, -36.171, -36.171, -36.171, -36.171, -36.171, -36.172, -36.172, 
    -36.172, -36.172, -36.172, -36.172, -36.172, -36.172, -36.172, -36.172, 
    -36.172, -36.173, -36.173, -36.173, -36.173, -36.173, -36.173, -36.173, 
    -36.173, -36.173, -36.174, -36.174, -36.174, -36.174, -36.174, -36.174, 
    -36.174, -36.174, -36.175, -36.175, -36.175, -36.175, -36.175, -36.175, 
    -36.176, -36.176, -36.176, -36.176, -36.176, -36.177, -36.177, -36.177, 
    -36.177, -36.178, -36.178, -36.179, -36.179, -36.18, -36.183, -36.185, 
    -36.186, -36.187, -36.188, -36.188, -36.189, -36.189, -36.19, -36.19, 
    -36.191, -36.192, -36.192, -36.193, -36.193, -36.194, -36.195, -36.195, 
    -36.196, -36.197, -36.197, -36.198, -36.199, -36.199, -36.2, -36.201, 
    -36.201, -36.202, -36.203, -36.204, -36.205, -36.206, -36.208, -36.21, 
    -36.211, -36.212, -36.212, -36.213, -36.213, -36.213, -36.214, -36.214, 
    -36.214, -36.215, -36.215, -36.215, -36.215, -36.216, -36.216, -36.216, 
    -36.216, -36.217, -36.217, -36.217, -36.217, -36.217, -36.218, -36.218, 
    -36.218, -36.218, -36.218, -36.219, -36.219, -36.219, -36.219, -36.219, 
    -36.219, -36.22, -36.22, -36.22, -36.22, -36.22, -36.221, -36.221, 
    -36.221, -36.221, -36.221, -36.221, -36.222, -36.222, -36.222, -36.222, 
    -36.222, -36.223, -36.223, -36.223, -36.223, -36.223, -36.224, -36.224, 
    -36.224, -36.224, -36.224, -36.225, -36.225, -36.225, -36.225, -36.225, 
    -36.226, -36.226, -36.226, -36.226, -36.227, -36.227, -36.227, -36.227, 
    -36.228, -36.228, -36.228, -36.229, -36.229, -36.229, -36.23, -36.23, 
    -36.23, -36.23, -36.231, -36.231, -36.231, -36.232, -36.232, -36.232, 
    -36.232, -36.233, -36.233, -36.233, -36.234, -36.234, -36.234, -36.234, 
    -36.234, -36.235, -36.235, -36.235, -36.235, -36.236, -36.236, -36.236, 
    -36.236, -36.236, -36.237, -36.237, -36.237, -36.237, -36.237, -36.237, 
    -36.238, -36.238, -36.238, -36.238, -36.238, -36.238, -36.239, -36.239, 
    -36.239, -36.239, -36.239, -36.239, -36.24, -36.24, -36.24, -36.24, 
    -36.24, -36.24, -36.24, -36.241, -36.241, -36.241, -36.241, -36.241, 
    -36.241, -36.242, -36.242, -36.242, -36.242, -36.242, -36.242, -36.242, 
    -36.243, -36.243, -36.243, -36.243, -36.243, -36.243, -36.243, -36.244, 
    -36.244, -36.244, -36.244, -36.244, -36.244, -36.245, -36.245, -36.245, 
    -36.245, -36.245, -36.245, -36.246, -36.246, -36.246, -36.246, -36.246, 
    -36.246, -36.247, -36.247, -36.247, -36.247, -36.247, -36.248, -36.248, 
    -36.248, -36.248, -36.248, -36.249, -36.249, -36.249, -36.249, -36.25, 
    -36.25, -36.25, -36.25, -36.251, -36.251, -36.251, -36.252, -36.252, 
    -36.252, -36.253, -36.253, -36.253, -36.254, -36.254, -36.254, -36.255, 
    -36.255, -36.255, -36.256, -36.256, -36.256, -36.257, -36.257, -36.257, 
    -36.257, -36.258, -36.258, -36.258, -36.258, -36.259, -36.259, -36.259, 
    -36.259, -36.26, -36.26, -36.26, -36.26, -36.26, -36.261, -36.261, 
    -36.261, -36.261, -36.261, -36.262, -36.262, -36.262, -36.262, -36.262, 
    -36.263, -36.263, -36.263, -36.263, -36.263, -36.264, -36.264, -36.264, 
    -36.264, -36.264, -36.265, -36.265, -36.265, -36.265, -36.265, -36.266, 
    -36.266, -36.266, -36.266, -36.266, -36.267, -36.267, -36.267, -36.267, 
    -36.267, -36.268, -36.268, -36.268, -36.268, -36.269, -36.269, -36.269, 
    -36.269, -36.269, -36.27, -36.27, -36.27, -36.27, -36.271, -36.271, 
    -36.271, -36.271, -36.272, -36.272, -36.272, -36.272, -36.273, -36.273, 
    -36.273, -36.273, -36.274, -36.274, -36.274, -36.274, -36.275, -36.275, 
    -36.275, -36.276, -36.276, -36.276, -36.276, -36.277, -36.277, -36.277, 
    -36.277, -36.278, -36.278, -36.278, -36.278, -36.279, -36.279, -36.279, 
    -36.279, -36.279, -36.28, -36.28, -36.28, -36.28, -36.281, -36.281, 
    -36.281, -36.281, -36.281, -36.282, -36.282, -36.282, -36.282, -36.282, 
    -36.282, -36.283, -36.283, -36.283, -36.283, -36.283, -36.284, -36.284, 
    -36.284, -36.284, -36.284, -36.284, -36.285, -36.285, -36.285, -36.285, 
    -36.285, -36.285, -36.286, -36.286, -36.286, -36.286, -36.286, -36.286, 
    -36.286, -36.287, -36.287, -36.287, -36.287, -36.287, -36.287, -36.288, 
    -36.288, -36.288, -36.288, -36.288, -36.288, -36.289, -36.289, -36.289, 
    -36.289, -36.289, -36.289, -36.29, -36.29, -36.29, -36.29, -36.29, 
    -36.29, -36.29, -36.291, -36.291, -36.291, -36.291, -36.291, -36.291, 
    -36.292, -36.292, -36.292, -36.292, -36.292, -36.292, -36.293, -36.293, 
    -36.293, -36.293, -36.293, -36.294, -36.294, -36.294, -36.294, -36.294, 
    -36.294, -36.295, -36.295, -36.295, -36.295, -36.295, -36.296, -36.296, 
    -36.296, -36.296, -36.296, -36.296, -36.297, -36.297, -36.297, -36.297, 
    -36.297, -36.298, -36.298, -36.298, -36.298, -36.298, -36.299, -36.299, 
    -36.299, -36.299, -36.3, -36.3, -36.3, -36.3, -36.3, -36.301, -36.301, 
    -36.301, -36.301, -36.301, -36.302, -36.302, -36.302, -36.302, -36.303, 
    -36.303, -36.303, -36.303, -36.303, -36.304, -36.304, -36.304, -36.304, 
    -36.305, -36.305, -36.305, -36.305, -36.305, -36.306, -36.306, -36.306, 
    -36.306, -36.307, -36.307, -36.307, -36.307, -36.307, -36.308, -36.308, 
    -36.308, -36.308, -36.308, -36.309, -36.309, -36.309, -36.309, -36.309, 
    -36.31, -36.31, -36.31, -36.31, -36.311, -36.311, -36.311, -36.311, 
    -36.311, -36.312, -36.312, -36.312, -36.312, -36.313, -36.313, -36.313, 
    -36.313, -36.313, -36.314, -36.314, -36.314, -36.314, -36.315, -36.315, 
    -36.315, -36.315, -36.316, -36.316, -36.316, -36.317, -36.317, -36.317, 
    -36.317, -36.318, -36.318, -36.318, -36.319, -36.319, -36.319, -36.319, 
    -36.32, -36.32, -36.32, -36.321, -36.321, -36.321, -36.322, -36.322, 
    -36.322, -36.323, -36.323, -36.323, -36.324, -36.324, -36.324, -36.324, 
    -36.325, -36.325, -36.325, -36.326, -36.326, -36.326, -36.326, -36.327, 
    -36.327, -36.327, -36.328, -36.328, -36.328, -36.328, -36.329, -36.329, 
    -36.329, -36.329, -36.33, -36.33, -36.33, -36.33, -36.331, -36.331, 
    -36.331, -36.331, -36.332, -36.332, -36.332, -36.332, -36.332, -36.333, 
    -36.333, -36.333, -36.333, -36.334, -36.334, -36.334, -36.334, -36.335, 
    -36.335, -36.335, -36.335, -36.335, -36.336, -36.336, -36.336, -36.336, 
    -36.336, -36.337, -36.337, -36.337, -36.337, -36.338, -36.338, -36.338, 
    -36.338, -36.338, -36.339, -36.339, -36.339, -36.339, -36.339, -36.34, 
    -36.34, -36.34, -36.34, -36.341, -36.341, -36.341, -36.341, -36.341, 
    -36.342, -36.342, -36.342, -36.342, -36.342, -36.343, -36.343, -36.343, 
    -36.343, -36.343, -36.344, -36.344, -36.344, -36.344, -36.344, -36.345, 
    -36.345, -36.345, -36.345, -36.345, -36.346, -36.346, -36.346, -36.346, 
    -36.346, -36.347, -36.347, -36.347, -36.347, -36.347, -36.348, -36.348, 
    -36.348, -36.348, -36.348, -36.348, -36.349, -36.349, -36.349, -36.349, 
    -36.349, -36.349, -36.35, -36.35, -36.35, -36.35, -36.35, -36.35, 
    -36.351, -36.351, -36.351, -36.351, -36.351, -36.351, -36.352, -36.352, 
    -36.352, -36.352, -36.352, -36.352, -36.353, -36.353, -36.353, -36.353, 
    -36.353, -36.353, -36.353, -36.354, -36.354, -36.354, -36.354, -36.354, 
    -36.354, -36.355, -36.355, -36.355, -36.355, -36.355, -36.355, -36.356, 
    -36.356, -36.356, -36.356, -36.356, -36.356, -36.356, -36.357, -36.357, 
    -36.357, -36.357, -36.357, -36.357, -36.358, -36.358, -36.358, -36.358, 
    -36.358, -36.358, -36.359, -36.359, -36.359, -36.359, -36.359, -36.359, 
    -36.36, -36.36, -36.36, -36.36, -36.36, -36.36, -36.361, -36.361, 
    -36.361, -36.361, -36.361, -36.361, -36.362, -36.362, -36.362, -36.362, 
    -36.362, -36.363, -36.363, -36.363, -36.363, -36.363, -36.364, -36.364, 
    -36.364, -36.364, -36.364, -36.364, -36.365, -36.365, -36.365, -36.365, 
    -36.365, -36.366, -36.366, -36.366, -36.366, -36.366, -36.367, -36.367, 
    -36.367, -36.367, -36.367, -36.368, -36.368, -36.368, -36.368, -36.368, 
    -36.369, -36.369, -36.369, -36.369, -36.369, -36.37, -36.37, -36.37, 
    -36.37, -36.371, -36.371, -36.371, -36.371, -36.371, -36.372, -36.372, 
    -36.372, -36.372, -36.372, -36.373, -36.373, -36.373, -36.373, -36.373, 
    -36.374, -36.374, -36.374, -36.374, -36.374, -36.374, -36.375, -36.375, 
    -36.375, -36.375, -36.375, -36.376, -36.376, -36.376, -36.376, -36.376, 
    -36.377, -36.377, -36.377, -36.377, -36.377, -36.377, -36.378, -36.378, 
    -36.378, -36.378, -36.378, -36.378, -36.379, -36.379, -36.379, -36.379, 
    -36.379, -36.379, -36.38, -36.38, -36.38, -36.38, -36.38, -36.38, 
    -36.381, -36.381, -36.381, -36.381, -36.381, -36.381, -36.382, -36.382, 
    -36.382, -36.382, -36.382, -36.382, -36.382, -36.383, -36.383, -36.383, 
    -36.383, -36.383, -36.383, -36.384, -36.384, -36.384, -36.384, -36.384, 
    -36.384, -36.385, -36.385, -36.385, -36.385, -36.385, -36.385, -36.386, 
    -36.386, -36.386, -36.386, -36.386, -36.387, -36.387, -36.387, -36.387, 
    -36.387, -36.387, -36.388, -36.388, -36.388, -36.388, -36.388, -36.388, 
    -36.389, -36.389, -36.389, -36.389, -36.389, -36.39, -36.39, -36.39, 
    -36.39, -36.39, -36.391, -36.391, -36.391, -36.391, -36.391, -36.392, 
    -36.392, -36.392, -36.392, -36.393, -36.393, -36.393, -36.393, -36.393, 
    -36.394, -36.394, -36.394, -36.394, -36.395, -36.395, -36.395, -36.395, 
    -36.395, -36.396, -36.396, -36.396, -36.396, -36.397, -36.397, -36.397, 
    -36.397, -36.398, -36.398, -36.398, -36.398, -36.399, -36.399, -36.399, 
    -36.399, -36.399, -36.4, -36.4, -36.4, -36.4, -36.401, -36.401, -36.401, 
    -36.401, -36.401, -36.402, -36.402, -36.402, -36.402, -36.402, -36.403, 
    -36.403, -36.403, -36.403, -36.403, -36.404, -36.404, -36.404, -36.404, 
    -36.404, -36.405, -36.405, -36.405, -36.405, -36.405, -36.405, -36.406, 
    -36.406, -36.406, -36.406, -36.406, -36.407, -36.407, -36.407, -36.407, 
    -36.407, -36.407, -36.408, -36.408, -36.408, -36.408, -36.408, -36.408, 
    -36.409, -36.409, -36.409, -36.409, -36.409, -36.41, -36.41, -36.41, 
    -36.41, -36.41, -36.41, -36.411, -36.411, -36.411, -36.411, -36.411, 
    -36.411, -36.412, -36.412, -36.412, -36.412, -36.412, -36.413, -36.413, 
    -36.413, -36.413, -36.413, -36.413, -36.414, -36.414, -36.414, -36.414, 
    -36.414, -36.415, -36.415, -36.415, -36.415, -36.415, -36.415, -36.416, 
    -36.416, -36.416, -36.416, -36.416, -36.417, -36.417, -36.417, -36.417, 
    -36.417, -36.417, -36.418, -36.418, -36.418, -36.418, -36.418, -36.419, 
    -36.419, -36.419, -36.419, -36.419, -36.419, -36.42, -36.42, -36.42, 
    -36.42, -36.42, -36.42, -36.421, -36.421, -36.421, -36.421, -36.421, 
    -36.421, -36.422, -36.422, -36.422, -36.422, -36.422, -36.422, -36.423, 
    -36.423, -36.423, -36.423, -36.423, -36.423, -36.423, -36.424, -36.424, 
    -36.424, -36.424, -36.424, -36.424, -36.424, -36.425, -36.425, -36.425, 
    -36.425, -36.425, -36.425, -36.425, -36.426, -36.426, -36.426, -36.426, 
    -36.426, -36.426, -36.426, -36.427, -36.427, -36.427, -36.427, -36.427, 
    -36.427, -36.427, -36.427, -36.428, -36.428, -36.428, -36.428, -36.428, 
    -36.428, -36.428, -36.429, -36.429, -36.429, -36.429, -36.429, -36.429, 
    -36.429, -36.43, -36.43, -36.43, -36.43, -36.43, -36.43, -36.43, -36.43, 
    -36.431, -36.431, -36.431, -36.431, -36.431, -36.431, -36.431, -36.432, 
    -36.432, -36.432, -36.432, -36.432, -36.432, -36.432, -36.433, -36.433, 
    -36.433, -36.433, -36.433, -36.433, -36.433, -36.434, -36.434, -36.434, 
    -36.434, -36.434, -36.434, -36.435, -36.435, -36.435, -36.435, -36.435, 
    -36.435, -36.436, -36.436, -36.436, -36.436, -36.436, -36.437, -36.437, 
    -36.437, -36.437, -36.437, -36.437, -36.438, -36.438, -36.438, -36.438, 
    -36.439, -36.439, -36.439, -36.439, -36.439, -36.44, -36.44, -36.44, 
    -36.44, -36.441, -36.441, -36.441, -36.441, -36.442, -36.442, -36.442, 
    -36.442, -36.442, -36.443, -36.443, -36.443, -36.443, -36.444, -36.444, 
    -36.444, -36.444, -36.445, -36.445, -36.445, -36.445, -36.445, -36.446, 
    -36.446, -36.446, -36.446, -36.446, -36.447, -36.447, -36.447, -36.447, 
    -36.448, -36.448, -36.448, -36.448, -36.448, -36.448, -36.449, -36.449, 
    -36.449, -36.449, -36.449, -36.45, -36.45, -36.45, -36.45, -36.45, 
    -36.451, -36.451, -36.451, -36.451, -36.451, -36.452, -36.452, -36.452, 
    -36.452, -36.452, -36.452, -36.453, -36.453, -36.453, -36.453, -36.453, 
    -36.454, -36.454, -36.454, -36.454, -36.454, -36.455, -36.455, -36.455, 
    -36.455, -36.455, -36.456, -36.456, -36.456, -36.456, -36.456, -36.457, 
    -36.457, -36.457, -36.457, -36.457, -36.457, -36.458, -36.458, -36.458, 
    -36.458, -36.458, -36.459, -36.459, -36.459, -36.459, -36.459, -36.46, 
    -36.46, -36.46, -36.46, -36.46, -36.461, -36.461, -36.461, -36.461, 
    -36.461, -36.462, -36.462, -36.462, -36.462, -36.462, -36.463, -36.463, 
    -36.463, -36.463, -36.463, -36.464, -36.464, -36.464, -36.464, -36.464, 
    -36.464, -36.465, -36.465, -36.465, -36.465, -36.465, -36.466, -36.466, 
    -36.466, -36.466, -36.466, -36.466, -36.467, -36.467, -36.467, -36.467, 
    -36.467, -36.468, -36.468, -36.468, -36.468, -36.468, -36.468, -36.469, 
    -36.469, -36.469, -36.469, -36.469, -36.47, -36.47, -36.47, -36.47, 
    -36.47, -36.47, -36.471, -36.471, -36.471, -36.471, -36.471, -36.471, 
    -36.472, -36.472, -36.472, -36.472, -36.472, -36.472, -36.473, -36.473, 
    -36.473, -36.473, -36.473, -36.473, -36.474, -36.474, -36.474, -36.474, 
    -36.474, -36.474, -36.475, -36.475, -36.475, -36.475, -36.475, -36.475, 
    -36.476, -36.476, -36.476, -36.476, -36.476, -36.476, -36.477, -36.477, 
    -36.477, -36.477, -36.477, -36.477, -36.478, -36.478, -36.478, -36.478, 
    -36.478, -36.478, -36.479, -36.479, -36.479, -36.479, -36.479, -36.479, 
    -36.48, -36.48, -36.48, -36.48, -36.48, -36.48, -36.481, -36.481, 
    -36.481, -36.481, -36.481, -36.481, -36.482, -36.482, -36.482, -36.482, 
    -36.482, -36.482, -36.483, -36.483, -36.483, -36.483, -36.483, -36.483, 
    -36.484, -36.484, -36.484, -36.484, -36.484, -36.484, -36.485, -36.485, 
    -36.485, -36.485, -36.485, -36.485, -36.486, -36.486, -36.486, -36.486, 
    -36.486, -36.486, -36.487, -36.487, -36.487, -36.487, -36.487, -36.487, 
    -36.488, -36.488, -36.488, -36.488, -36.488, -36.489, -36.489, -36.489, 
    -36.489, -36.489, -36.489, -36.49, -36.49, -36.49, -36.49, -36.49, 
    -36.49, -36.491, -36.491, -36.491, -36.491, -36.491, -36.491, -36.492, 
    -36.492, -36.492, -36.492, -36.492, -36.492, -36.493, -36.493, -36.493, 
    -36.493, -36.493, -36.493, -36.493, -36.494, -36.494, -36.494, -36.494, 
    -36.494, -36.494, -36.495, -36.495, -36.495, -36.495, -36.495, -36.495, 
    -36.495, -36.496, -36.496, -36.496, -36.496, -36.496, -36.496, -36.497, 
    -36.497, -36.497, -36.497, -36.497, -36.497, -36.497, -36.498, -36.498, 
    -36.498, -36.498, -36.498, -36.498, -36.498, -36.499, -36.499, -36.499, 
    -36.499, -36.499, -36.499, -36.499, -36.5, -36.5, -36.5, -36.5, -36.5, 
    -36.5, -36.5, -36.501, -36.501, -36.501, -36.501, -36.501, -36.501, 
    -36.501, -36.502, -36.502, -36.502, -36.502, -36.502, -36.502, -36.502, 
    -36.503, -36.503, -36.503, -36.503, -36.503, -36.503, -36.503, -36.504, 
    -36.504, -36.504, -36.504, -36.504, -36.504, -36.504, -36.505, -36.505, 
    -36.505, -36.505, -36.505, -36.505, -36.505, -36.506, -36.506, -36.506, 
    -36.506, -36.506, -36.506, -36.506, -36.507, -36.507, -36.507, -36.507, 
    -36.507, -36.507, -36.507, -36.508, -36.508, -36.508, -36.508, -36.508, 
    -36.508, -36.508, -36.509, -36.509, -36.509, -36.509, -36.509, -36.509, 
    -36.51, -36.51, -36.51, -36.51, -36.51, -36.51, -36.511, -36.511, 
    -36.511, -36.511, -36.511, -36.511, -36.512, -36.512, -36.512, -36.512, 
    -36.512, -36.512, -36.513, -36.513, -36.513, -36.513, -36.513, -36.513, 
    -36.514, -36.514, -36.514, -36.514, -36.514, -36.514, -36.515, -36.515, 
    -36.515, -36.515, -36.515, -36.516, -36.516, -36.516, -36.516, -36.516, 
    -36.516, -36.517, -36.517, -36.517, -36.517, -36.517, -36.518, -36.518, 
    -36.518, -36.518, -36.518, -36.519, -36.519, -36.519, -36.519, -36.519, 
    -36.52, -36.52, -36.52, -36.52, -36.52, -36.521, -36.521, -36.521, 
    -36.521, -36.521, -36.521, -36.522, -36.522, -36.522, -36.522, -36.522, 
    -36.523, -36.523, -36.523, -36.523, -36.523, -36.523, -36.524, -36.524, 
    -36.524, -36.524, -36.524, -36.524, -36.525, -36.525, -36.525, -36.525, 
    -36.525, -36.525, -36.526, -36.526, -36.526, -36.526, -36.526, -36.526, 
    -36.526, -36.527, -36.527, -36.527, -36.527, -36.527, -36.527, -36.527, 
    -36.528, -36.528, -36.528, -36.528, -36.528, -36.528, -36.529, -36.529, 
    -36.529, -36.529, -36.529, -36.529, -36.529, -36.53, -36.53, -36.53, 
    -36.53, -36.53, -36.53, -36.53, -36.531, -36.531, -36.531, -36.531, 
    -36.531, -36.531, -36.531, -36.532, -36.532, -36.532, -36.532, -36.532, 
    -36.532, -36.532, -36.532, -36.533, -36.533, -36.533, -36.533, -36.533, 
    -36.533, -36.533, -36.534, -36.534, -36.534, -36.534, -36.534, -36.534, 
    -36.534, -36.535, -36.535, -36.535, -36.535, -36.535, -36.535, -36.535, 
    -36.536, -36.536, -36.536, -36.536, -36.536, -36.536, -36.536, -36.537, 
    -36.537, -36.537, -36.537, -36.537, -36.537, -36.537, -36.537, -36.538, 
    -36.538, -36.538, -36.538, -36.538, -36.538, -36.538, -36.539, -36.539, 
    -36.539, -36.539, -36.539, -36.539, -36.539, -36.54, -36.54, -36.54, 
    -36.54, -36.54, -36.54, -36.54, -36.54, -36.541, -36.541, -36.541, 
    -36.541, -36.541, -36.541, -36.541, -36.542, -36.542, -36.542, -36.542, 
    -36.542, -36.542, -36.542, -36.542, -36.543, -36.543, -36.543, -36.543, 
    -36.543, -36.543, -36.543, -36.543, -36.544, -36.544, -36.544, -36.544, 
    -36.544, -36.544, -36.544, -36.545, -36.545, -36.545, -36.545, -36.545, 
    -36.545, -36.545, -36.545, -36.546, -36.546, -36.546, -36.546, -36.546, 
    -36.546, -36.546, -36.546, -36.547, -36.547, -36.547, -36.547, -36.547, 
    -36.547, -36.547, -36.548, -36.548, -36.548, -36.548, -36.548, -36.548, 
    -36.548, -36.548, -36.549, -36.549, -36.549, -36.549, -36.549, -36.549, 
    -36.549, -36.549, -36.55, -36.55, -36.55, -36.55, -36.55, -36.55, -36.55, 
    -36.551, -36.551, -36.551, -36.551, -36.551, -36.551, -36.551, -36.552, 
    -36.552, -36.552, -36.552, -36.552, -36.552, -36.552, -36.553, -36.553, 
    -36.553, -36.553, -36.553, -36.553, -36.553, -36.554, -36.554, -36.554, 
    -36.554, -36.554, -36.554, -36.554, -36.555, -36.555, -36.555, -36.555, 
    -36.555, -36.555, -36.556, -36.556, -36.556, -36.556, -36.556, -36.556, 
    -36.556, -36.557, -36.557, -36.557, -36.557, -36.557, -36.557, -36.558, 
    -36.558, -36.558, -36.558, -36.558, -36.558, -36.559, -36.559, -36.559, 
    -36.559, -36.559, -36.559, -36.56, -36.56, -36.56, -36.56, -36.56, 
    -36.56, -36.561, -36.561, -36.561, -36.561, -36.561, -36.561, -36.562, 
    -36.562, -36.562, -36.562, -36.562, -36.562, -36.563, -36.563, -36.563, 
    -36.563, -36.563, -36.563, -36.564, -36.564, -36.564, -36.564, -36.564, 
    -36.564, -36.564, -36.565, -36.565, -36.565, -36.565, -36.565, -36.565, 
    -36.566, -36.566, -36.566, -36.566, -36.566, -36.566, -36.567, -36.567, 
    -36.567, -36.567, -36.567, -36.567, -36.567, -36.568, -36.568, -36.568, 
    -36.568, -36.568, -36.568, -36.568, -36.569, -36.569, -36.569, -36.569, 
    -36.569, -36.569, -36.569, -36.57, -36.57, -36.57, -36.57, -36.57, 
    -36.57, -36.57, -36.571, -36.571, -36.571, -36.571, -36.571, -36.571, 
    -36.571, -36.571, -36.572, -36.572, -36.572, -36.572, -36.572, -36.572, 
    -36.572, -36.572, -36.573, -36.573, -36.573, -36.573, -36.573, -36.573, 
    -36.573, -36.573, -36.574, -36.574, -36.574, -36.574, -36.574, -36.574, 
    -36.574, -36.574, -36.574, -36.575, -36.575, -36.575, -36.575, -36.575, 
    -36.575, -36.575, -36.575, -36.575, -36.576, -36.576, -36.576, -36.576, 
    -36.576, -36.576, -36.576, -36.576, -36.576, -36.577, -36.577, -36.577, 
    -36.577, -36.577, -36.577, -36.577, -36.577, -36.577, -36.577, -36.578, 
    -36.578, -36.578, -36.578, -36.578, -36.578, -36.578, -36.578, -36.578, 
    -36.578, -36.579, -36.579, -36.579, -36.579, -36.579, -36.579, -36.579, 
    -36.579, -36.579, -36.579, -36.58, -36.58, -36.58, -36.58, -36.58, 
    -36.58, -36.58, -36.58, -36.58, -36.58, -36.58, -36.581, -36.581, 
    -36.581, -36.581, -36.581, -36.581, -36.581, -36.581, -36.581, -36.581, 
    -36.581, -36.582, -36.582, -36.582, -36.582, -36.582, -36.582, -36.582, 
    -36.582, -36.582, -36.582, -36.583, -36.583, -36.583, -36.583, -36.583, 
    -36.583, -36.583, -36.583, -36.583, -36.583, -36.583, -36.584, -36.584, 
    -36.584, -36.584, -36.584, -36.584, -36.584, -36.584, -36.584, -36.584, 
    -36.584, -36.585, -36.585, -36.585, -36.585, -36.585, -36.585, -36.585, 
    -36.585, -36.585, -36.585, -36.585, -36.586, -36.586, -36.586, -36.586, 
    -36.586, -36.586, -36.586, -36.586, -36.586, -36.586, -36.586, -36.586, 
    -36.587, -36.587, -36.587, -36.587, -36.587, -36.587, -36.587, -36.587, 
    -36.587, -36.587, -36.588, -36.588, -36.588, -36.588, -36.588, -36.588, 
    -36.588, -36.588, -36.588, -36.588, -36.588, -36.589, -36.589, -36.589, 
    -36.589, -36.589, -36.589, -36.589, -36.589, -36.589, -36.589, -36.589, 
    -36.59, -36.59, -36.59, -36.59, -36.59, -36.59, -36.59, -36.59, -36.59, 
    -36.59, -36.59, -36.591, -36.591, -36.591, -36.591, -36.591, -36.591, 
    -36.591, -36.591, -36.591, -36.591, -36.592, -36.592, -36.592, -36.592, 
    -36.592, -36.592, -36.592, -36.592, -36.592, -36.592, -36.593, -36.593, 
    -36.593, -36.593, -36.593, -36.593, -36.593, -36.593, -36.593, -36.593, 
    -36.594, -36.594, -36.594, -36.594, -36.594, -36.594, -36.594, -36.594, 
    -36.594, -36.595, -36.595, -36.595, -36.595, -36.595, -36.595, -36.595, 
    -36.595, -36.595, -36.596, -36.596, -36.596, -36.596, -36.596, -36.596, 
    -36.596, -36.596, -36.596, -36.597, -36.597, -36.597, -36.597, -36.597, 
    -36.597, -36.597, -36.597, -36.598, -36.598, -36.598, -36.598, -36.598, 
    -36.598, -36.598, -36.598, -36.599, -36.599, -36.599, -36.599, -36.599, 
    -36.599, -36.599, -36.6, -36.6, -36.6, -36.6, -36.6, -36.6, -36.601, 
    -36.601, -36.601, -36.601, -36.601, -36.601, -36.602, -36.602, -36.602, 
    -36.602, -36.602, -36.603, -36.603, -36.603, -36.603, -36.603, -36.604, 
    -36.604, -36.604, -36.604, -36.605, -36.605, -36.605, -36.606, -36.606, 
    -36.606, -36.606, -36.607, -36.607, -36.607, -36.608, -36.608, -36.608, 
    -36.609, -36.609, -36.609, -36.61, -36.61, -36.61, -36.611, -36.611, 
    -36.612, -36.612, -36.612, -36.613, -36.613, -36.613, -36.614, -36.614, 
    -36.614, -36.615, -36.615, -36.616, -36.616, -36.616, -36.617, -36.617, 
    -36.617, -36.617, -36.618, -36.618, -36.618, -36.619, -36.619, -36.619, 
    -36.619, -36.62, -36.62, -36.62, -36.62, -36.62, -36.621, -36.621, 
    -36.621, -36.621, -36.622, -36.622, -36.622, -36.622, -36.622, -36.622, 
    -36.623, -36.623, -36.623, -36.623, -36.623, -36.623, -36.624, -36.624, 
    -36.624, -36.624, -36.624, -36.624, -36.625, -36.625, -36.625, -36.625, 
    -36.625, -36.625, -36.626, -36.626, -36.626, -36.626, -36.626, -36.626, 
    -36.626, -36.627, -36.627, -36.627, -36.627, -36.627, -36.627, -36.627, 
    -36.628, -36.628, -36.628, -36.628, -36.628, -36.628, -36.628, -36.629, 
    -36.629, -36.629, -36.629, -36.629, -36.629, -36.629, -36.63, -36.63, 
    -36.63, -36.63, -36.63, -36.63, -36.63, -36.631, -36.631, -36.631, 
    -36.631, -36.631, -36.631, -36.631, -36.632, -36.632, -36.632, -36.632, 
    -36.632, -36.632, -36.632, -36.632, -36.633, -36.633, -36.633, -36.633, 
    -36.633, -36.633, -36.633, -36.634, -36.634, -36.634, -36.634, -36.634, 
    -36.634, -36.634, -36.635, -36.635, -36.635, -36.635, -36.635, -36.635, 
    -36.635, -36.635, -36.636, -36.636, -36.636, -36.636, -36.636, -36.636, 
    -36.636, -36.637, -36.637, -36.637, -36.637, -36.637, -36.637, -36.637, 
    -36.637, -36.638, -36.638, -36.638, -36.638, -36.638, -36.638, -36.638, 
    -36.639, -36.639, -36.639, -36.639, -36.639, -36.639, -36.639, -36.639, 
    -36.64, -36.64, -36.64, -36.64, -36.64, -36.64, -36.64, -36.64, -36.641, 
    -36.641, -36.641, -36.641, -36.641, -36.641, -36.641, -36.642, -36.642, 
    -36.642, -36.642, -36.642, -36.642, -36.642, -36.642, -36.643, -36.643, 
    -36.643, -36.643, -36.643, -36.643, -36.643, -36.644, -36.644, -36.644, 
    -36.644, -36.644, -36.644, -36.644, -36.645, -36.645, -36.645, -36.645, 
    -36.645, -36.645, -36.645, -36.646, -36.646, -36.646, -36.646, -36.646, 
    -36.646, -36.647, -36.647, -36.647, -36.647, -36.647, -36.647, -36.648, 
    -36.648, -36.648, -36.648, -36.648, -36.648, -36.649, -36.649, -36.649, 
    -36.649, -36.649, -36.65, -36.65, -36.65, -36.65, -36.65, -36.651, 
    -36.651, -36.651, -36.651, -36.651, -36.652, -36.652, -36.652, -36.652, 
    -36.653, -36.653, -36.653, -36.653, -36.654, -36.654, -36.654, -36.654, 
    -36.655, -36.655, -36.655, -36.655, -36.655, -36.656, -36.656, -36.656, 
    -36.656, -36.657, -36.657, -36.657, -36.657, -36.658, -36.658, -36.658, 
    -36.658, -36.658, -36.659, -36.659, -36.659, -36.659, -36.659, -36.66, 
    -36.66, -36.66, -36.66, -36.661, -36.661, -36.661, -36.661, -36.661, 
    -36.662, -36.662, -36.662, -36.662, -36.662, -36.663, -36.663, -36.663, 
    -36.663, -36.664, -36.664, -36.664, -36.664, -36.664, -36.665, -36.665, 
    -36.665, -36.665, -36.666, -36.666, -36.666, -36.666, -36.667, -36.667, 
    -36.667, -36.667, -36.667, -36.668, -36.668, -36.668, -36.668, -36.669, 
    -36.669, -36.669, -36.669, -36.67, -36.67, -36.67, -36.67, -36.671, 
    -36.671, -36.671, -36.671, -36.672, -36.672, -36.672, -36.672, -36.673, 
    -36.673, -36.673, -36.673, -36.673, -36.674, -36.674, -36.674, -36.674, 
    -36.675, -36.675, -36.675, -36.675, -36.675, -36.676, -36.676, -36.676, 
    -36.676, -36.677, -36.677, -36.677, -36.677, -36.677, -36.678, -36.678, 
    -36.678, -36.678, -36.678, -36.679, -36.679, -36.679, -36.679, -36.679, 
    -36.68, -36.68, -36.68, -36.68, -36.681, -36.681, -36.681, -36.681, 
    -36.681, -36.682, -36.682, -36.682, -36.682, -36.683, -36.683, -36.683, 
    -36.683, -36.683, -36.684, -36.684, -36.684, -36.684, -36.685, -36.685, 
    -36.685, -36.685, -36.685, -36.686, -36.686, -36.686, -36.686, -36.686, 
    -36.687, -36.687, -36.687, -36.687, -36.687, -36.688, -36.688, -36.688, 
    -36.688, -36.688, -36.689, -36.689, -36.689, -36.689, -36.689, -36.69, 
    -36.69, -36.69, -36.69, -36.69, -36.691, -36.691, -36.691, -36.691, 
    -36.691, -36.691, -36.692, -36.692, -36.692, -36.692, -36.692, -36.692, 
    -36.693, -36.693, -36.693, -36.693, -36.693, -36.693, -36.694, -36.694, 
    -36.694, -36.694, -36.694, -36.695, -36.695, -36.695, -36.695, -36.695, 
    -36.695, -36.696, -36.696, -36.696, -36.696, -36.696, -36.696, -36.697, 
    -36.697, -36.697, -36.697, -36.697, -36.697, -36.698, -36.698, -36.698, 
    -36.698, -36.698, -36.698, -36.699, -36.699, -36.699, -36.699, -36.699, 
    -36.699, -36.7, -36.7, -36.7, -36.7, -36.7, -36.7, -36.701, -36.701, 
    -36.701, -36.701, -36.701, -36.701, -36.702, -36.702, -36.702, -36.702, 
    -36.702, -36.702, -36.703, -36.703, -36.703, -36.703, -36.703, -36.704, 
    -36.704, -36.704, -36.704, -36.704, -36.705, -36.705, -36.705, -36.705, 
    -36.705, -36.706, -36.706, -36.706, -36.706, -36.706, -36.707, -36.707, 
    -36.707, -36.707, -36.707, -36.708, -36.708, -36.708, -36.708, -36.709, 
    -36.709, -36.709, -36.709, -36.71, -36.71, -36.71, -36.71, -36.711, 
    -36.711, -36.711, -36.711, -36.711, -36.712, -36.712, -36.712, -36.712, 
    -36.713, -36.713, -36.713, -36.713, -36.713, -36.714, -36.714, -36.714, 
    -36.714, -36.714, -36.715, -36.715, -36.715, -36.715, -36.715, -36.716, 
    -36.716, -36.716, -36.716, -36.716, -36.716, -36.717, -36.717, -36.717, 
    -36.717, -36.717, -36.718, -36.718, -36.718, -36.718, -36.718, -36.718, 
    -36.719, -36.719, -36.719, -36.719, -36.719, -36.719, -36.719, -36.72, 
    -36.72, -36.72, -36.72, -36.72, -36.72, -36.721, -36.721, -36.721, 
    -36.721, -36.721, -36.721, -36.721, -36.722, -36.722, -36.722, -36.722, 
    -36.722, -36.722, -36.723, -36.723, -36.723, -36.723, -36.723, -36.723, 
    -36.723, -36.724, -36.724, -36.724, -36.724, -36.724, -36.724, -36.725, 
    -36.725, -36.725, -36.725, -36.725, -36.725, -36.725, -36.726, -36.726, 
    -36.726, -36.726, -36.726, -36.726, -36.727, -36.727, -36.728, -36.728, 
    -36.729, -36.729, -36.73, -36.73, -36.731, -36.732, -36.732, -36.733, 
    -36.733, -36.734, -36.734, -36.735, -36.735, -36.736, -36.737, -36.737, 
    -36.738, -36.738, -36.739, -36.739, -36.74, -36.74, -36.741, -36.742, 
    -36.742, -36.743, -36.743, -36.744, -36.745, -36.745, -36.746, -36.746, 
    -36.747, -36.747, -36.748, -36.749, -36.749, -36.75, -36.75, -36.751, 
    -36.751, -36.752, -36.753, -36.753, -36.754, -36.754, -36.755, -36.755, 
    -36.756, -36.756, -36.757, -36.758, -36.758, -36.759, -36.759, -36.76, 
    -36.76, -36.761, -36.762, -36.762, -36.763, -36.763, -36.764, -36.764, 
    -36.765, -36.766, -36.766, -36.767, -36.767, -36.768, -36.769, -36.769, 
    -36.77, -36.77, -36.771, -36.771, -36.772, -36.773, -36.773, -36.774, 
    -36.774, -36.775, -36.775, -36.776, -36.777, -36.777, -36.778, -36.778, 
    -36.779, -36.779, -36.78, -36.781, -36.781, -36.782, -36.782, -36.783, 
    -36.783, -36.784, -36.785, -36.785, -36.786, -36.786, -36.787, -36.788, 
    -36.788, -36.789, -36.789, -36.79, -36.79, -36.791, -36.792, -36.792, 
    -36.793, -36.793, -36.794, -36.795, -36.795, -36.796, -36.796, -36.797, 
    -36.797, -36.798, -36.799, -36.799, -36.8, -36.8, -36.801, -36.802, 
    -36.802, -36.803, -36.803, -36.804, -36.804, -36.805, -36.806, -36.806, 
    -36.807, -36.807, -36.808, -36.808, -36.809, -36.81, -36.81, -36.811, 
    -36.811, -36.812, -36.813, -36.813, -36.814, -36.814, -36.815, -36.816, 
    -36.816, -36.817, -36.817, -36.818, -36.819, -36.819, -36.82, -36.82, 
    -36.821, -36.822, -36.822, -36.823, -36.823, -36.824, -36.825, -36.825, 
    -36.826, -36.826, -36.827, -36.828, -36.828, -36.829, -36.829, -36.83, 
    -36.831, -36.831, -36.832, -36.832, -36.833, -36.834, -36.834, -36.835, 
    -36.835, -36.836, -36.837, -36.837, -36.838, -36.838, -36.839, -36.84, 
    -36.84, -36.841, -36.842, -36.842, -36.843, -36.843, -36.844, -36.845, 
    -36.845, -36.846, -36.846, -36.847, -36.848, -36.848, -36.849, -36.849, 
    -36.85, -36.851, -36.851, -36.852, -36.853, -36.853, -36.854, -36.855, 
    -36.855, -36.856, -36.856, -36.857, -36.858, -36.858, -36.859, -36.86, 
    -36.86, -36.861, -36.862, -36.862, -36.863, -36.864, -36.864, -36.865, 
    -36.866, -36.866, -36.867, -36.868, -36.868, -36.869, -36.869, -36.87, 
    -36.871, -36.871, -36.872, -36.873, -36.873, -36.874, -36.875, -36.875, 
    -36.876, -36.877, -36.877, -36.878, -36.878, -36.879, -36.88, -36.88, 
    -36.881, -36.882, -36.882, -36.883, -36.883, -36.884, -36.885, -36.885, 
    -36.886, -36.887, -36.887, -36.888, -36.888, -36.889, -36.89, -36.89, 
    -36.891, -36.891, -36.892, -36.893, -36.893, -36.894, -36.894, -36.895, 
    -36.896, -36.896, -36.897, -36.897, -36.898, -36.899, -36.899, -36.9, 
    -36.9, -36.901, -36.902, -36.902, -36.903, -36.903, -36.904, -36.905, 
    -36.905, -36.906, -36.907, -36.907, -36.908, -36.908, -36.909, -36.91, 
    -36.91, -36.911, -36.911, -36.912, -36.913, -36.913, -36.914, -36.915, 
    -36.915, -36.916, -36.917, -36.917, -36.918, -36.919, -36.919, -36.92, 
    -36.92, -36.921, -36.922, -36.922, -36.923, -36.924, -36.924, -36.925, 
    -36.926, -36.926, -36.927, -36.928, -36.928, -36.929, -36.93, -36.93, 
    -36.931, -36.932, -36.932, -36.933, -36.934, -36.935, -36.935, -36.936, 
    -36.937, -36.937, -36.938, -36.939, -36.939, -36.94, -36.941, -36.941, 
    -36.942, -36.943, -36.943, -36.944, -36.944, -36.945, -36.946, -36.946, 
    -36.947, -36.948, -36.948, -36.949, -36.95, -36.95, -36.951, -36.952, 
    -36.952, -36.953, -36.954, -36.954, -36.955, -36.956, -36.956, -36.957, 
    -36.958, -36.958, -36.959, -36.959, -36.96, -36.961, -36.961, -36.962, 
    -36.963, -36.963, -36.964, -36.965, -36.965, -36.966, -36.967, -36.967, 
    -36.968, -36.968, -36.969, -36.97, -36.97, -36.971, -36.972, -36.972, 
    -36.973, -36.974, -36.974, -36.975, -36.976, -36.976, -36.977, -36.978, 
    -36.978, -36.979, -36.98, -36.98, -36.981, -36.982, -36.982, -36.983, 
    -36.984, -36.984, -36.985, -36.986, -36.986, -36.987, -36.988, -36.988, 
    -36.989, -36.99, -36.99, -36.991, -36.992, -36.992, -36.993, -36.994, 
    -36.994, -36.995, -36.996, -36.996, -36.997, -36.998, -36.998, -36.999, 
    -37, -37, -37.001, -37.002, -37.002, -37.003, -37.004, -37.004, -37.005, 
    -37.006, -37.006, -37.007, -37.008, -37.008, -37.009, -37.01, -37.01, 
    -37.011, -37.012, -37.012, -37.013, -37.014, -37.014, -37.015, -37.016, 
    -37.016, -37.017, -37.018, -37.019, -37.019, -37.02, -37.021, -37.021, 
    -37.022, -37.023, -37.024, -37.024, -37.025, -37.026, -37.026, -37.027, 
    -37.028, -37.028, -37.029, -37.03, -37.031, -37.031, -37.032, -37.033, 
    -37.033, -37.034, -37.035, -37.035, -37.036, -37.037, -37.038, -37.038, 
    -37.039, -37.04, -37.04, -37.041, -37.042, -37.042, -37.043, -37.044, 
    -37.044, -37.045, -37.046, -37.046, -37.047, -37.048, -37.048, -37.049, 
    -37.05, -37.05, -37.051, -37.052, -37.052, -37.053, -37.054, -37.055, 
    -37.055, -37.056, -37.057, -37.057, -37.058, -37.059, -37.06, -37.06, 
    -37.061, -37.062, -37.062, -37.063, -37.064, -37.065, -37.065, -37.066, 
    -37.067, -37.068, -37.068, -37.069, -37.07, -37.07, -37.071, -37.072, 
    -37.073, -37.073, -37.074, -37.075, -37.075, -37.076, -37.077, -37.078, 
    -37.078, -37.079, -37.08, -37.081, -37.081, -37.082, -37.083, -37.083, 
    -37.084, -37.085, -37.086, -37.086, -37.087, -37.088, -37.088, -37.089, 
    -37.09, -37.091, -37.091, -37.092, -37.093, -37.093, -37.094, -37.095, 
    -37.096, -37.096, -37.097, -37.098, -37.098, -37.099, -37.1, -37.1, 
    -37.101, -37.102, -37.103, -37.103, -37.104, -37.105, -37.105, -37.106, 
    -37.107, -37.108, -37.108, -37.109, -37.11, -37.11, -37.111, -37.112, 
    -37.113, -37.113, -37.114, -37.115, -37.116, -37.116, -37.117, -37.118, 
    -37.119, -37.119, -37.12, -37.121, -37.122, -37.122, -37.123, -37.124, 
    -37.125, -37.125, -37.126, -37.127, -37.128, -37.128, -37.129, -37.13, 
    -37.131, -37.131, -37.132, -37.133, -37.134, -37.134, -37.135, -37.136, 
    -37.137, -37.137, -37.138, -37.139, -37.14, -37.14, -37.141, -37.142, 
    -37.143, -37.143, -37.144, -37.145, -37.146, -37.146, -37.147, -37.148, 
    -37.149, -37.149, -37.15, -37.151, -37.152, -37.152, -37.153, -37.154, 
    -37.155, -37.155, -37.156, -37.157, -37.157, -37.158, -37.159, -37.16, 
    -37.16, -37.161, -37.162, -37.163, -37.163, -37.164, -37.165, -37.166, 
    -37.166, -37.167, -37.168, -37.169, -37.169, -37.17, -37.171, -37.171, 
    -37.172, -37.173, -37.174, -37.174, -37.175, -37.176, -37.177, -37.177, 
    -37.178, -37.179, -37.18, -37.181, -37.181, -37.182, -37.183, -37.184, 
    -37.184, -37.185, -37.186, -37.187, -37.188, -37.188, -37.189, -37.19, 
    -37.191, -37.191, -37.192, -37.193, -37.194, -37.195, -37.195, -37.196, 
    -37.197, -37.198, -37.199, -37.199, -37.2, -37.201, -37.202, -37.202, 
    -37.203, -37.204, -37.205, -37.206, -37.206, -37.207, -37.208, -37.209, 
    -37.209, -37.21, -37.211, -37.212, -37.212, -37.213, -37.214, -37.215, 
    -37.216, -37.216, -37.217, -37.218, -37.219, -37.219, -37.22, -37.221, 
    -37.222, -37.223, -37.223, -37.224, -37.225, -37.226, -37.226, -37.227, 
    -37.228, -37.229, -37.229, -37.23, -37.231, -37.232, -37.233, -37.233, 
    -37.234, -37.235, -37.236, -37.236, -37.237, -37.238, -37.239, -37.239, 
    -37.24, -37.241, -37.242, -37.243, -37.243, -37.244, -37.245, -37.246, 
    -37.246, -37.247, -37.248, -37.249, -37.249, -37.25, -37.251, -37.252, 
    -37.253, -37.253, -37.254, -37.255, -37.256, -37.256, -37.257, -37.258, 
    -37.259, -37.26, -37.26, -37.261, -37.262, -37.263, -37.264, -37.264, 
    -37.265, -37.266, -37.267, -37.268, -37.268, -37.269, -37.27, -37.271, 
    -37.272, -37.272, -37.273, -37.274, -37.275, -37.275, -37.276, -37.277, 
    -37.278, -37.279, -37.279, -37.28, -37.281, -37.282, -37.283, -37.283, 
    -37.284, -37.285, -37.286, -37.287, -37.287, -37.288, -37.289, -37.29, 
    -37.291, -37.291, -37.292, -37.293, -37.294, -37.295, -37.295, -37.296, 
    -37.297, -37.298, -37.299, -37.299, -37.3, -37.301, -37.302, -37.303, 
    -37.303, -37.304, -37.305, -37.306, -37.307, -37.307, -37.308, -37.309, 
    -37.31, -37.311, -37.311, -37.312, -37.313, -37.314, -37.315, -37.315, 
    -37.316, -37.317, -37.318, -37.319, -37.319, -37.32, -37.321, -37.322, 
    -37.323, -37.324, -37.324, -37.325, -37.326, -37.327, -37.328, -37.328, 
    -37.329, -37.33, -37.331, -37.332, -37.332, -37.333, -37.334, -37.335, 
    -37.336, -37.336, -37.337, -37.338, -37.339, -37.34, -37.34, -37.341, 
    -37.342, -37.343, -37.344, -37.345, -37.345, -37.346, -37.347, -37.348, 
    -37.349, -37.349, -37.35, -37.351, -37.352, -37.353, -37.353, -37.354, 
    -37.355, -37.356, -37.357, -37.357, -37.358, -37.359, -37.36, -37.361, 
    -37.361, -37.362, -37.363, -37.364, -37.365, -37.365, -37.366, -37.367, 
    -37.368, -37.369, -37.369, -37.37, -37.371, -37.372, -37.373, -37.374, 
    -37.374, -37.375, -37.376, -37.377, -37.378, -37.378, -37.379, -37.38, 
    -37.381, -37.382, -37.383, -37.383, -37.384, -37.385, -37.386, -37.387, 
    -37.387, -37.388, -37.389, -37.39, -37.391, -37.391, -37.392, -37.393, 
    -37.394, -37.395, -37.396, -37.396, -37.397, -37.398, -37.399, -37.4, 
    -37.4, -37.401, -37.402, -37.403, -37.404, -37.405, -37.405, -37.406, 
    -37.407, -37.408, -37.409, -37.409, -37.41, -37.411, -37.412, -37.413, 
    -37.414, -37.414, -37.415, -37.416, -37.417, -37.418, -37.418, -37.419, 
    -37.42, -37.421, -37.422, -37.422, -37.423, -37.424, -37.425, -37.426, 
    -37.427, -37.427, -37.428, -37.429, -37.43, -37.431, -37.431, -37.432, 
    -37.433, -37.434, -37.435, -37.435, -37.436, -37.437, -37.438, -37.439, 
    -37.44, -37.44, -37.441, -37.442, -37.443, -37.444, -37.444, -37.445, 
    -37.446, -37.447, -37.448, -37.449, -37.449, -37.45, -37.451, -37.452, 
    -37.453, -37.454, -37.454, -37.455, -37.456, -37.457, -37.458, -37.459, 
    -37.459, -37.46, -37.461, -37.462, -37.463, -37.464, -37.464, -37.465, 
    -37.466, -37.467, -37.468, -37.468, -37.469, -37.47, -37.471, -37.472, 
    -37.473, -37.473, -37.474, -37.475, -37.476, -37.477, -37.478, -37.478, 
    -37.479, -37.48, -37.481, -37.482, -37.482, -37.483, -37.484, -37.485, 
    -37.486, -37.487, -37.487, -37.488, -37.489, -37.49, -37.491, -37.491, 
    -37.492, -37.493, -37.494, -37.495, -37.496, -37.496, -37.497, -37.498, 
    -37.499, -37.5, -37.501, -37.501, -37.502, -37.503, -37.504, -37.505, 
    -37.505, -37.506, -37.507, -37.508, -37.509, -37.51, -37.51, -37.511, 
    -37.512, -37.513, -37.514, -37.515, -37.515, -37.516, -37.517, -37.518, 
    -37.519, -37.52, -37.52, -37.521, -37.522, -37.523, -37.524, -37.524, 
    -37.525, -37.526, -37.527, -37.528, -37.529, -37.529, -37.53, -37.531, 
    -37.532, -37.533, -37.534, -37.534, -37.535, -37.536, -37.537, -37.538, 
    -37.539, -37.539, -37.54, -37.541, -37.542, -37.543, -37.544, -37.544, 
    -37.545, -37.546, -37.547, -37.548, -37.548, -37.549, -37.55, -37.551, 
    -37.552, -37.553, -37.553, -37.554, -37.555, -37.556, -37.557, -37.558, 
    -37.558, -37.559, -37.56, -37.561, -37.562, -37.563, -37.563, -37.564, 
    -37.565, -37.566, -37.567, -37.568, -37.568, -37.569, -37.57, -37.571, 
    -37.572, -37.573, -37.573, -37.574, -37.575, -37.576, -37.577, -37.578, 
    -37.578, -37.579, -37.58, -37.581, -37.582, -37.583, -37.583, -37.584, 
    -37.585, -37.586, -37.587, -37.588, -37.588, -37.589, -37.59, -37.591, 
    -37.592, -37.593, -37.594, -37.594, -37.595, -37.596, -37.597, -37.598, 
    -37.599, -37.599, -37.6, -37.601, -37.602, -37.603, -37.604, -37.604, 
    -37.605, -37.606, -37.607, -37.608, -37.609, -37.609, -37.61, -37.611, 
    -37.612, -37.613, -37.613, -37.614, -37.615, -37.616, -37.617, -37.618, 
    -37.618, -37.619, -37.62, -37.621, -37.622, -37.622, -37.623, -37.624, 
    -37.625, -37.626, -37.627, -37.627, -37.628, -37.629, -37.63, -37.631, 
    -37.632, -37.633, -37.633, -37.634, -37.635, -37.636, -37.637, -37.638, 
    -37.638, -37.639, -37.64, -37.641, -37.642, -37.643, -37.643, -37.644, 
    -37.645, -37.646, -37.647, -37.648, -37.648, -37.649, -37.65, -37.651, 
    -37.652, -37.653, -37.653, -37.654, -37.655, -37.656, -37.657, -37.658, 
    -37.658, -37.659, -37.66, -37.661, -37.662, -37.663, -37.663, -37.664, 
    -37.665, -37.666, -37.667, -37.667, -37.668, -37.669, -37.67, -37.671, 
    -37.672, -37.672, -37.673, -37.674, -37.675, -37.676, -37.677, -37.677, 
    -37.678, -37.679, -37.68, -37.681, -37.682, -37.682, -37.683, -37.684, 
    -37.685, -37.686, -37.687, -37.687, -37.688, -37.689, -37.69, -37.691, 
    -37.692, -37.693, -37.693, -37.694, -37.695, -37.696, -37.697, -37.698, 
    -37.698, -37.699, -37.7, -37.701, -37.702, -37.703, -37.704, -37.704, 
    -37.705, -37.706, -37.707, -37.708, -37.709, -37.709, -37.71, -37.711, 
    -37.712, -37.713, -37.714, -37.714, -37.715, -37.716, -37.717, -37.718, 
    -37.719, -37.719, -37.72, -37.721, -37.722, -37.723, -37.724, -37.724, 
    -37.725, -37.726, -37.727, -37.728, -37.729, -37.729, -37.73, -37.731, 
    -37.732, -37.733, -37.734, -37.734, -37.735, -37.736, -37.737, -37.738, 
    -37.739, -37.739, -37.74, -37.741, -37.742, -37.743, -37.744, -37.744, 
    -37.745, -37.746, -37.747, -37.748, -37.749, -37.749, -37.75, -37.751, 
    -37.752, -37.753, -37.754, -37.754, -37.755, -37.756, -37.757, -37.758, 
    -37.759, -37.759, -37.76, -37.761, -37.762, -37.763, -37.763, -37.764, 
    -37.765, -37.766, -37.767, -37.768, -37.768, -37.769, -37.77, -37.771, 
    -37.772, -37.773, -37.773, -37.774, -37.775, -37.776, -37.777, -37.778, 
    -37.778, -37.779, -37.78, -37.781, -37.782, -37.783, -37.784, -37.784, 
    -37.785, -37.786, -37.787, -37.788, -37.789, -37.789, -37.79, -37.791, 
    -37.792, -37.793, -37.794, -37.794, -37.795, -37.796, -37.797, -37.798, 
    -37.799, -37.799, -37.8, -37.801, -37.802, -37.803, -37.804, -37.804, 
    -37.805, -37.806, -37.807, -37.808, -37.809, -37.809, -37.81, -37.811, 
    -37.812, -37.813, -37.814, -37.815, -37.815, -37.816, -37.817, -37.818, 
    -37.819, -37.82, -37.82, -37.821, -37.822, -37.823, -37.824, -37.825, 
    -37.825, -37.826, -37.827, -37.828, -37.829, -37.83, -37.83, -37.831, 
    -37.832, -37.833, -37.834, -37.835, -37.835, -37.836, -37.837, -37.838, 
    -37.839, -37.84, -37.84, -37.841, -37.842, -37.843, -37.844, -37.845, 
    -37.846, -37.846, -37.847, -37.848, -37.849, -37.85, -37.851, -37.851, 
    -37.852, -37.853, -37.854, -37.855, -37.856, -37.856, -37.857, -37.858, 
    -37.859, -37.86, -37.861, -37.861, -37.862, -37.863, -37.864, -37.865, 
    -37.866, -37.867, -37.867, -37.868, -37.869, -37.87, -37.871, -37.872, 
    -37.872, -37.873, -37.874, -37.875, -37.876, -37.877, -37.878, -37.878, 
    -37.879, -37.88, -37.881, -37.882, -37.883, -37.883, -37.884, -37.885, 
    -37.886, -37.887, -37.888, -37.888, -37.889, -37.89, -37.891, -37.892, 
    -37.893, -37.893, -37.894, -37.895, -37.896, -37.897, -37.898, -37.898, 
    -37.899, -37.9, -37.901, -37.902, -37.903, -37.903, -37.904, -37.905, 
    -37.906, -37.907, -37.908, -37.909, -37.909, -37.91, -37.911, -37.912, 
    -37.913, -37.914, -37.914, -37.915, -37.916, -37.917, -37.918, -37.919, 
    -37.919, -37.92, -37.921, -37.922, -37.923, -37.924, -37.924, -37.925, 
    -37.926, -37.927, -37.928, -37.929 ;

 azimuth_tp =
  136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 
    136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.54, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 
    136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 136.56, 
    136.56, 136.56, 136.56, 136.55, 136.55, 136.55, 136.55, 136.55, 136.55, 
    136.55, 136.55, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 136.59, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 
    136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.6, 136.61, 
    136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 
    136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 
    136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 
    136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 136.61, 
    136.61, 136.61, 136.61, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 136.62, 
    136.62, 136.62, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 136.63, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 
    136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.64, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 136.65, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 136.66, 
    136.66, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 
    136.67, 136.67, 136.67, 136.67, 136.67, 136.67, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 136.68, 
    136.68, 136.68, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 
    136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.69, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 
    136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.7, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 136.71, 
    136.71, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 136.72, 
    136.72, 136.72, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 136.73, 
    136.73, 136.73, 136.73, 136.73, 136.73, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 136.74, 
    136.74, 136.74, 136.74, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 136.75, 
    136.75, 136.75, 136.75, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 136.76, 
    136.76, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 
    136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.77, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 
    136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.78, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 136.79, 
    136.79, 136.79, 136.79, 136.79, 136.79, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 136.8, 
    136.8, 136.8, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 
    136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 
    136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 
    136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 
    136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 
    136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.81, 136.82, 
    136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 
    136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 
    136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 
    136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 
    136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.82, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 136.83, 
    136.83, 136.83, 136.83, 136.83, 136.84, 136.84, 136.84, 136.84, 136.84, 
    136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 
    136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 
    136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 
    136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 136.84, 
    136.84, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 
    136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 
    136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 
    136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 
    136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 136.85, 
    136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 
    136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 
    136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 
    136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 
    136.86, 136.86, 136.86, 136.86, 136.86, 136.86, 136.87, 136.87, 136.87, 
    136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 
    136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 
    136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 
    136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.87, 136.88, 
    136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 
    136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 
    136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 
    136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 136.88, 
    136.88, 136.88, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 
    136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 
    136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 
    136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 136.89, 
    136.89, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 
    136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 
    136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 
    136.9, 136.9, 136.9, 136.9, 136.9, 136.9, 136.91, 136.91, 136.91, 136.91, 
    136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 
    136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 
    136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 136.91, 
    136.91, 136.91, 136.91, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 
    136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 
    136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 
    136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.92, 136.93, 
    136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 
    136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 
    136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 136.93, 
    136.93, 136.93, 136.93, 136.93, 136.93, 136.94, 136.94, 136.94, 136.94, 
    136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 
    136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 
    136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.94, 136.95, 
    136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 
    136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 
    136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 136.95, 
    136.95, 136.95, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 
    136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 
    136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 136.96, 
    136.96, 136.96, 136.96, 136.96, 136.96, 136.97, 136.97, 136.97, 136.97, 
    136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 
    136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 
    136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.97, 136.98, 
    136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 
    136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 
    136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 136.98, 
    136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 
    136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 
    136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 136.99, 
    136.99, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 
    137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 
    137, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 
    137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 
    137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 137.01, 
    137.01, 137.01, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 
    137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 
    137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 137.02, 
    137.02, 137.02, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 
    137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 
    137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 137.03, 
    137.03, 137.03, 137.03, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 
    137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 
    137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 137.04, 
    137.04, 137.04, 137.04, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 
    137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 
    137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 137.05, 
    137.05, 137.05, 137.05, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 
    137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 
    137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 137.06, 
    137.06, 137.06, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 
    137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 
    137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 137.07, 
    137.07, 137.07, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 
    137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 
    137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 137.08, 
    137.08, 137.08, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 
    137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 
    137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 137.09, 
    137.09, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 
    137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 
    137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.1, 137.11, 137.11, 
    137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 
    137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 
    137.11, 137.11, 137.11, 137.11, 137.11, 137.11, 137.12, 137.12, 137.12, 
    137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 
    137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 137.12, 
    137.12, 137.12, 137.12, 137.12, 137.12, 137.13, 137.13, 137.13, 137.13, 
    137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 
    137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 137.13, 
    137.13, 137.13, 137.13, 137.13, 137.14, 137.14, 137.14, 137.14, 137.14, 
    137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 
    137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 137.14, 
    137.14, 137.14, 137.14, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 
    137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 
    137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 137.15, 
    137.15, 137.15, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 
    137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 
    137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 137.16, 
    137.16, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 
    137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 
    137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 137.17, 
    137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 
    137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 
    137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.18, 137.19, 
    137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 
    137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 
    137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.19, 137.2, 137.2, 
    137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 
    137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 137.2, 
    137.2, 137.2, 137.2, 137.2, 137.21, 137.21, 137.21, 137.21, 137.21, 
    137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 
    137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 137.21, 
    137.21, 137.21, 137.21, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 
    137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 
    137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 137.22, 
    137.22, 137.22, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 
    137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 
    137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 137.23, 
    137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 
    137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 
    137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.24, 137.25, 
    137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 
    137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 
    137.25, 137.25, 137.25, 137.25, 137.25, 137.25, 137.26, 137.26, 137.26, 
    137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 
    137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 137.26, 
    137.26, 137.26, 137.26, 137.26, 137.26, 137.27, 137.27, 137.27, 137.27, 
    137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 
    137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 137.27, 
    137.27, 137.27, 137.27, 137.27, 137.28, 137.28, 137.28, 137.28, 137.28 ;

 impact_L1 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 impact_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 impact =
  6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3976e+06, 
    6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 
    6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 6.3977e+06, 
    6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 
    6.3977e+06, 6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 
    6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 
    6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 
    6.398e+06, 6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 
    6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 
    6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 
    6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 
    6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3984e+06, 
    6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 
    6.3984e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3986e+06, 6.3986e+06, 
    6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 
    6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 
    6.3987e+06, 6.3987e+06, 6.3988e+06, 6.3988e+06, 6.3988e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 
    6.3989e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 
    6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 
    6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3993e+06, 
    6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 
    6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 
    6.3994e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 
    6.3995e+06, 6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 
    6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3998e+06, 
    6.3998e+06, 6.3998e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 
    6.3999e+06, 6.3999e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4e+06, 6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 
    6.4001e+06, 6.4001e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4002e+06, 6.4002e+06, 6.4002e+06, 6.4002e+06, 6.4003e+06, 6.4003e+06, 
    6.4003e+06, 6.4003e+06, 6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 
    6.4004e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 6.4005e+06, 
    6.4005e+06, 6.4005e+06, 6.4006e+06, 6.4006e+06, 6.4006e+06, 6.4006e+06, 
    6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 
    6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4009e+06, 
    6.4009e+06, 6.4009e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 
    6.401e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 6.4011e+06, 6.4011e+06, 
    6.4011e+06, 6.4011e+06, 6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4012e+06, 
    6.4012e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4013e+06, 6.4013e+06, 6.4013e+06, 6.4014e+06, 6.4014e+06, 6.4014e+06, 
    6.4014e+06, 6.4014e+06, 6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 
    6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 
    6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4017e+06, 
    6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 
    6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 
    6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 
    6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4022e+06, 6.4022e+06, 6.4022e+06, 6.4023e+06, 6.4023e+06, 
    6.4023e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4024e+06, 6.4024e+06, 
    6.4024e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 
    6.4027e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 6.4028e+06, 
    6.4028e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 
    6.403e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4031e+06, 6.4031e+06, 6.4031e+06, 6.4032e+06, 6.4032e+06, 
    6.4032e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4033e+06, 
    6.4033e+06, 6.4033e+06, 6.4034e+06, 6.4034e+06, 6.4034e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 
    6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 
    6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4038e+06, 
    6.4038e+06, 6.4038e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 
    6.4039e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 6.404e+06, 6.404e+06, 
    6.404e+06, 6.404e+06, 6.4041e+06, 6.4041e+06, 6.4041e+06, 6.4041e+06, 
    6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4043e+06, 6.4043e+06, 6.4043e+06, 6.4043e+06, 6.4044e+06, 6.4044e+06, 
    6.4044e+06, 6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4045e+06, 
    6.4045e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4048e+06, 
    6.4048e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 6.4049e+06, 
    6.4049e+06, 6.4049e+06, 6.405e+06, 6.405e+06, 6.405e+06, 6.405e+06, 
    6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 
    6.4052e+06, 6.4052e+06, 6.4052e+06, 6.4053e+06, 6.4053e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 
    6.4055e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 6.4056e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 
    6.4058e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 6.4059e+06, 6.4059e+06, 
    6.4059e+06, 6.406e+06, 6.406e+06, 6.406e+06, 6.406e+06, 6.4061e+06, 
    6.4061e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 6.4062e+06, 
    6.4062e+06, 6.4062e+06, 6.4063e+06, 6.4063e+06, 6.4063e+06, 6.4063e+06, 
    6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 
    6.4065e+06, 6.4065e+06, 6.4065e+06, 6.4066e+06, 6.4066e+06, 6.4066e+06, 
    6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 
    6.4068e+06, 6.4068e+06, 6.4068e+06, 6.4069e+06, 6.4069e+06, 6.4069e+06, 
    6.407e+06, 6.407e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4071e+06, 6.4072e+06, 6.4072e+06, 6.4072e+06, 6.4072e+06, 6.4073e+06, 
    6.4073e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 
    6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4077e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4078e+06, 6.4078e+06, 6.4079e+06, 6.4079e+06, 6.4079e+06, 
    6.4079e+06, 6.408e+06, 6.408e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4081e+06, 6.4081e+06, 6.4081e+06, 6.4082e+06, 6.4082e+06, 6.4082e+06, 
    6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 
    6.4084e+06, 6.4084e+06, 6.4084e+06, 6.4085e+06, 6.4085e+06, 6.4085e+06, 
    6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4087e+06, 
    6.4087e+06, 6.4087e+06, 6.4088e+06, 6.4088e+06, 6.4088e+06, 6.4089e+06, 
    6.4089e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.409e+06, 
    6.4091e+06, 6.4091e+06, 6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4092e+06, 
    6.4092e+06, 6.4093e+06, 6.4093e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4094e+06, 6.4095e+06, 6.4095e+06, 6.4095e+06, 6.4095e+06, 6.4096e+06, 
    6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 6.4097e+06, 6.4098e+06, 
    6.4098e+06, 6.4098e+06, 6.4098e+06, 6.4099e+06, 6.4099e+06, 6.4099e+06, 
    6.41e+06, 6.41e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4102e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 
    6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 6.4104e+06, 6.4105e+06, 
    6.4105e+06, 6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4106e+06, 
    6.4107e+06, 6.4107e+06, 6.4107e+06, 6.4107e+06, 6.4108e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 
    6.411e+06, 6.411e+06, 6.4111e+06, 6.4111e+06, 6.4111e+06, 6.4111e+06, 
    6.4112e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4113e+06, 6.4113e+06, 
    6.4114e+06, 6.4114e+06, 6.4114e+06, 6.4115e+06, 6.4115e+06, 6.4115e+06, 
    6.4116e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4118e+06, 6.4118e+06, 6.4119e+06, 6.4119e+06, 6.4119e+06, 
    6.412e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 6.4121e+06, 6.4121e+06, 
    6.4122e+06, 6.4122e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4123e+06, 
    6.4124e+06, 6.4124e+06, 6.4124e+06, 6.4124e+06, 6.4125e+06, 6.4125e+06, 
    6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4127e+06, 
    6.4127e+06, 6.4128e+06, 6.4128e+06, 6.4128e+06, 6.4129e+06, 6.4129e+06, 
    6.4129e+06, 6.413e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4132e+06, 6.4132e+06, 6.4132e+06, 6.4133e+06, 
    6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 6.4134e+06, 6.4135e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 
    6.4137e+06, 6.4137e+06, 6.4138e+06, 6.4138e+06, 6.4138e+06, 6.4139e+06, 
    6.4139e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.414e+06, 
    6.4141e+06, 6.4141e+06, 6.4141e+06, 6.4142e+06, 6.4142e+06, 6.4142e+06, 
    6.4143e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4146e+06, 
    6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 6.4148e+06, 6.4148e+06, 
    6.4149e+06, 6.4149e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.415e+06, 
    6.4151e+06, 6.4151e+06, 6.4151e+06, 6.4152e+06, 6.4152e+06, 6.4152e+06, 
    6.4153e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4154e+06, 
    6.4155e+06, 6.4155e+06, 6.4155e+06, 6.4156e+06, 6.4156e+06, 6.4156e+06, 
    6.4157e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4158e+06, 6.4158e+06, 
    6.4159e+06, 6.4159e+06, 6.416e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 
    6.4161e+06, 6.4161e+06, 6.4162e+06, 6.4162e+06, 6.4162e+06, 6.4163e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 
    6.4165e+06, 6.4165e+06, 6.4166e+06, 6.4166e+06, 6.4166e+06, 6.4167e+06, 
    6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 
    6.4171e+06, 6.4172e+06, 6.4172e+06, 6.4172e+06, 6.4173e+06, 6.4173e+06, 
    6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4177e+06, 6.4177e+06, 
    6.4178e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 6.4179e+06, 6.418e+06, 
    6.418e+06, 6.418e+06, 6.4181e+06, 6.4181e+06, 6.4181e+06, 6.4182e+06, 
    6.4182e+06, 6.4182e+06, 6.4183e+06, 6.4183e+06, 6.4183e+06, 6.4184e+06, 
    6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4185e+06, 6.4186e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 
    6.4188e+06, 6.4189e+06, 6.4189e+06, 6.4189e+06, 6.419e+06, 6.419e+06, 
    6.419e+06, 6.4191e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4193e+06, 6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4194e+06, 
    6.4195e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 6.4196e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 
    6.4199e+06, 6.4199e+06, 6.42e+06, 6.42e+06, 6.42e+06, 6.4201e+06, 
    6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 6.4203e+06, 
    6.4203e+06, 6.4204e+06, 6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 
    6.4205e+06, 6.4206e+06, 6.4206e+06, 6.4206e+06, 6.4207e+06, 6.4207e+06, 
    6.4208e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.4209e+06, 6.4209e+06, 
    6.421e+06, 6.421e+06, 6.421e+06, 6.4211e+06, 6.4211e+06, 6.4212e+06, 
    6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4213e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 
    6.4216e+06, 6.4217e+06, 6.4217e+06, 6.4217e+06, 6.4218e+06, 6.4218e+06, 
    6.4218e+06, 6.4219e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.422e+06, 
    6.422e+06, 6.4221e+06, 6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4222e+06, 
    6.4223e+06, 6.4223e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 
    6.4227e+06, 6.4227e+06, 6.4228e+06, 6.4228e+06, 6.4228e+06, 6.4229e+06, 
    6.4229e+06, 6.423e+06, 6.423e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 
    6.4231e+06, 6.4232e+06, 6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4233e+06, 
    6.4234e+06, 6.4234e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 6.4236e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 
    6.4238e+06, 6.4238e+06, 6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 
    6.424e+06, 6.4241e+06, 6.4241e+06, 6.4241e+06, 6.4242e+06, 6.4242e+06, 
    6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4244e+06, 6.4244e+06, 
    6.4245e+06, 6.4245e+06, 6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4246e+06, 
    6.4247e+06, 6.4247e+06, 6.4248e+06, 6.4248e+06, 6.4248e+06, 6.4249e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 
    6.4251e+06, 6.4252e+06, 6.4252e+06, 6.4252e+06, 6.4253e+06, 6.4253e+06, 
    6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4256e+06, 6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4257e+06, 
    6.4258e+06, 6.4258e+06, 6.4259e+06, 6.4259e+06, 6.4259e+06, 6.426e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 
    6.4262e+06, 6.4263e+06, 6.4263e+06, 6.4263e+06, 6.4264e+06, 6.4264e+06, 
    6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 6.4266e+06, 6.4266e+06, 
    6.4267e+06, 6.4267e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4268e+06, 
    6.4269e+06, 6.4269e+06, 6.427e+06, 6.427e+06, 6.427e+06, 6.4271e+06, 
    6.4271e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4275e+06, 
    6.4275e+06, 6.4276e+06, 6.4276e+06, 6.4277e+06, 6.4277e+06, 6.4277e+06, 
    6.4278e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.428e+06, 6.4281e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 
    6.4282e+06, 6.4283e+06, 6.4283e+06, 6.4283e+06, 6.4284e+06, 6.4284e+06, 
    6.4284e+06, 6.4285e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4286e+06, 
    6.4287e+06, 6.4287e+06, 6.4287e+06, 6.4288e+06, 6.4288e+06, 6.4289e+06, 
    6.4289e+06, 6.4289e+06, 6.429e+06, 6.429e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 
    6.4293e+06, 6.4294e+06, 6.4294e+06, 6.4295e+06, 6.4295e+06, 6.4295e+06, 
    6.4296e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 6.4298e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.4299e+06, 6.4299e+06, 6.43e+06, 
    6.43e+06, 6.4301e+06, 6.4301e+06, 6.4301e+06, 6.4302e+06, 6.4302e+06, 
    6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4304e+06, 6.4305e+06, 6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4306e+06, 
    6.4307e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 6.4308e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 
    6.4311e+06, 6.4311e+06, 6.4312e+06, 6.4312e+06, 6.4313e+06, 6.4313e+06, 
    6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4317e+06, 
    6.4318e+06, 6.4318e+06, 6.4319e+06, 6.4319e+06, 6.4319e+06, 6.432e+06, 
    6.432e+06, 6.432e+06, 6.4321e+06, 6.4321e+06, 6.4322e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 
    6.4324e+06, 6.4325e+06, 6.4325e+06, 6.4326e+06, 6.4326e+06, 6.4326e+06, 
    6.4327e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.4329e+06, 6.433e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 
    6.4331e+06, 6.4331e+06, 6.4332e+06, 6.4332e+06, 6.4332e+06, 6.4333e+06, 
    6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4335e+06, 
    6.4335e+06, 6.4336e+06, 6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4337e+06, 
    6.4338e+06, 6.4338e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 6.434e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4342e+06, 
    6.4342e+06, 6.4343e+06, 6.4343e+06, 6.4343e+06, 6.4344e+06, 6.4344e+06, 
    6.4345e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 6.4346e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 
    6.4349e+06, 6.4349e+06, 6.435e+06, 6.435e+06, 6.435e+06, 6.4351e+06, 
    6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 6.4353e+06, 
    6.4353e+06, 6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4355e+06, 
    6.4356e+06, 6.4356e+06, 6.4356e+06, 6.4357e+06, 6.4357e+06, 6.4357e+06, 
    6.4358e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 
    6.436e+06, 6.436e+06, 6.4361e+06, 6.4361e+06, 6.4361e+06, 6.4362e+06, 
    6.4362e+06, 6.4363e+06, 6.4363e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4364e+06, 6.4365e+06, 6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4366e+06, 
    6.4367e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 6.4368e+06, 6.4368e+06, 
    6.4369e+06, 6.4369e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 
    6.4371e+06, 6.4371e+06, 6.4372e+06, 6.4372e+06, 6.4372e+06, 6.4373e+06, 
    6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 6.4375e+06, 6.4375e+06, 
    6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4377e+06, 
    6.4377e+06, 6.4378e+06, 6.4378e+06, 6.4379e+06, 6.4379e+06, 6.4379e+06, 
    6.438e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 6.4381e+06, 6.4382e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 
    6.4384e+06, 6.4385e+06, 6.4385e+06, 6.4385e+06, 6.4386e+06, 6.4386e+06, 
    6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.439e+06, 
    6.4391e+06, 6.4391e+06, 6.4392e+06, 6.4392e+06, 6.4392e+06, 6.4393e+06, 
    6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4394e+06, 6.4394e+06, 6.4395e+06, 
    6.4395e+06, 6.4396e+06, 6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4397e+06, 
    6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 6.4399e+06, 6.4399e+06, 
    6.44e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4401e+06, 
    6.4402e+06, 6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 
    6.4404e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 6.4406e+06, 6.4406e+06, 
    6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4408e+06, 
    6.4408e+06, 6.4409e+06, 6.4409e+06, 6.441e+06, 6.441e+06, 6.441e+06, 
    6.4411e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 6.4412e+06, 6.4413e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 
    6.4415e+06, 6.4416e+06, 6.4416e+06, 6.4416e+06, 6.4417e+06, 6.4417e+06, 
    6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.442e+06, 6.442e+06, 6.4421e+06, 6.4421e+06, 6.4421e+06, 
    6.4422e+06, 6.4422e+06, 6.4423e+06, 6.4423e+06, 6.4423e+06, 6.4424e+06, 
    6.4424e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4426e+06, 6.4427e+06, 6.4427e+06, 6.4427e+06, 6.4428e+06, 6.4428e+06, 
    6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 6.443e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4432e+06, 
    6.4433e+06, 6.4433e+06, 6.4434e+06, 6.4434e+06, 6.4434e+06, 6.4435e+06, 
    6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4437e+06, 6.4438e+06, 6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 
    6.4439e+06, 6.444e+06, 6.444e+06, 6.4441e+06, 6.4441e+06, 6.4441e+06, 
    6.4442e+06, 6.4442e+06, 6.4442e+06 ;

 impact_opt =
  6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3863e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3867e+06, 
    6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 6.3869e+06, 
    6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 
    6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 
    6.3874e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3883e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.3889e+06, 6.3889e+06, 6.3889e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 
    6.3896e+06, 6.3896e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 
    6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3906e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3908e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 
    6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 
    6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3928e+06, 6.3928e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3935e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 
    6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 
    6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.395e+06, 6.395e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 6.3951e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 6.3958e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.3959e+06, 6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.396e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 6.3962e+06, 
    6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3968e+06, 
    6.3968e+06, 6.3968e+06, 6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 
    6.3971e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 
    6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3972e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 6.3976e+06, 
    6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 
    6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 6.3977e+06, 
    6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 
    6.3977e+06, 6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 
    6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 
    6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 6.398e+06, 
    6.398e+06, 6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 
    6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 6.3981e+06, 
    6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3982e+06, 
    6.3982e+06, 6.3982e+06, 6.3982e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 
    6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3983e+06, 6.3984e+06, 
    6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 6.3984e+06, 
    6.3984e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3985e+06, 6.3986e+06, 6.3986e+06, 
    6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 6.3986e+06, 
    6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3987e+06, 
    6.3987e+06, 6.3987e+06, 6.3988e+06, 6.3988e+06, 6.3988e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 
    6.3989e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 
    6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3991e+06, 
    6.3991e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3993e+06, 
    6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 6.3993e+06, 
    6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 
    6.3994e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 
    6.3995e+06, 6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 
    6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3998e+06, 
    6.3998e+06, 6.3998e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 
    6.3999e+06, 6.3999e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4e+06, 6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 
    6.4001e+06, 6.4001e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4002e+06, 6.4002e+06, 6.4002e+06, 6.4002e+06, 6.4003e+06, 6.4003e+06, 
    6.4003e+06, 6.4003e+06, 6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 
    6.4004e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 6.4005e+06, 
    6.4005e+06, 6.4005e+06, 6.4006e+06, 6.4006e+06, 6.4006e+06, 6.4006e+06, 
    6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 6.4007e+06, 
    6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4008e+06, 6.4009e+06, 
    6.4009e+06, 6.4009e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 
    6.401e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 6.4011e+06, 6.4011e+06, 
    6.4011e+06, 6.4011e+06, 6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4012e+06, 
    6.4012e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4013e+06, 6.4013e+06, 6.4013e+06, 6.4014e+06, 6.4014e+06, 6.4014e+06, 
    6.4014e+06, 6.4014e+06, 6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 
    6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 
    6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4016e+06, 6.4017e+06, 
    6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 6.4017e+06, 
    6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 6.4018e+06, 
    6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 6.402e+06, 
    6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4022e+06, 6.4022e+06, 6.4022e+06, 6.4023e+06, 6.4023e+06, 
    6.4023e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4024e+06, 6.4024e+06, 
    6.4024e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 
    6.4027e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 6.4028e+06, 
    6.4028e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 6.4029e+06, 
    6.403e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4031e+06, 6.4031e+06, 6.4031e+06, 6.4032e+06, 6.4032e+06, 
    6.4032e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4033e+06, 
    6.4033e+06, 6.4033e+06, 6.4034e+06, 6.4034e+06, 6.4034e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 6.4035e+06, 
    6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 6.4036e+06, 
    6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4037e+06, 6.4038e+06, 
    6.4038e+06, 6.4038e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 
    6.4039e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 6.404e+06, 6.404e+06, 
    6.404e+06, 6.404e+06, 6.4041e+06, 6.4041e+06, 6.4041e+06, 6.4041e+06, 
    6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4043e+06, 6.4043e+06, 6.4043e+06, 6.4043e+06, 6.4044e+06, 6.4044e+06, 
    6.4044e+06, 6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4045e+06, 
    6.4045e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4047e+06, 6.4048e+06, 
    6.4048e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 6.4049e+06, 
    6.4049e+06, 6.4049e+06, 6.405e+06, 6.405e+06, 6.405e+06, 6.405e+06, 
    6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 
    6.4052e+06, 6.4052e+06, 6.4052e+06, 6.4053e+06, 6.4053e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 
    6.4055e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 6.4056e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 
    6.4058e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 6.4059e+06, 6.4059e+06, 
    6.4059e+06, 6.406e+06, 6.406e+06, 6.406e+06, 6.406e+06, 6.4061e+06, 
    6.4061e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 6.4062e+06, 
    6.4062e+06, 6.4062e+06, 6.4063e+06, 6.4063e+06, 6.4063e+06, 6.4063e+06, 
    6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 
    6.4065e+06, 6.4065e+06, 6.4065e+06, 6.4066e+06, 6.4066e+06, 6.4066e+06, 
    6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 
    6.4068e+06, 6.4068e+06, 6.4068e+06, 6.4069e+06, 6.4069e+06, 6.4069e+06, 
    6.407e+06, 6.407e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4071e+06, 6.4072e+06, 6.4072e+06, 6.4072e+06, 6.4072e+06, 6.4073e+06, 
    6.4073e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 
    6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4077e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4078e+06, 6.4078e+06, 6.4079e+06, 6.4079e+06, 6.4079e+06, 
    6.4079e+06, 6.408e+06, 6.408e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4081e+06, 6.4081e+06, 6.4081e+06, 6.4082e+06, 6.4082e+06, 6.4082e+06, 
    6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 
    6.4084e+06, 6.4084e+06, 6.4084e+06, 6.4085e+06, 6.4085e+06, 6.4085e+06, 
    6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4087e+06, 
    6.4087e+06, 6.4087e+06, 6.4088e+06, 6.4088e+06, 6.4088e+06, 6.4089e+06, 
    6.4089e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.409e+06, 
    6.4091e+06, 6.4091e+06, 6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4092e+06, 
    6.4092e+06, 6.4093e+06, 6.4093e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4094e+06, 6.4095e+06, 6.4095e+06, 6.4095e+06, 6.4095e+06, 6.4096e+06, 
    6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 6.4097e+06, 6.4098e+06, 
    6.4098e+06, 6.4098e+06, 6.4098e+06, 6.4099e+06, 6.4099e+06, 6.4099e+06, 
    6.41e+06, 6.41e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4102e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 
    6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 6.4104e+06, 6.4105e+06, 
    6.4105e+06, 6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4106e+06, 
    6.4107e+06, 6.4107e+06, 6.4107e+06, 6.4107e+06, 6.4108e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 
    6.411e+06, 6.411e+06, 6.4111e+06, 6.4111e+06, 6.4111e+06, 6.4111e+06, 
    6.4112e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4113e+06, 6.4113e+06, 
    6.4114e+06, 6.4114e+06, 6.4114e+06, 6.4115e+06, 6.4115e+06, 6.4115e+06, 
    6.4116e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4118e+06, 6.4118e+06, 6.4119e+06, 6.4119e+06, 6.4119e+06, 
    6.412e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 6.4121e+06, 6.4121e+06, 
    6.4122e+06, 6.4122e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4123e+06, 
    6.4124e+06, 6.4124e+06, 6.4124e+06, 6.4124e+06, 6.4125e+06, 6.4125e+06, 
    6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4127e+06, 
    6.4127e+06, 6.4128e+06, 6.4128e+06, 6.4128e+06, 6.4129e+06, 6.4129e+06, 
    6.4129e+06, 6.413e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4132e+06, 6.4132e+06, 6.4132e+06, 6.4133e+06, 
    6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 6.4134e+06, 6.4135e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 
    6.4137e+06, 6.4137e+06, 6.4138e+06, 6.4138e+06, 6.4138e+06, 6.4139e+06, 
    6.4139e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.414e+06, 
    6.4141e+06, 6.4141e+06, 6.4141e+06, 6.4142e+06, 6.4142e+06, 6.4142e+06, 
    6.4143e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4146e+06, 
    6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 6.4148e+06, 6.4148e+06, 
    6.4149e+06, 6.4149e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.415e+06, 
    6.4151e+06, 6.4151e+06, 6.4151e+06, 6.4152e+06, 6.4152e+06, 6.4152e+06, 
    6.4153e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4154e+06, 
    6.4155e+06, 6.4155e+06, 6.4155e+06, 6.4156e+06, 6.4156e+06, 6.4156e+06, 
    6.4157e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4158e+06, 6.4158e+06, 
    6.4159e+06, 6.4159e+06, 6.416e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 
    6.4161e+06, 6.4161e+06, 6.4162e+06, 6.4162e+06, 6.4162e+06, 6.4163e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 
    6.4165e+06, 6.4165e+06, 6.4166e+06, 6.4166e+06, 6.4166e+06, 6.4167e+06, 
    6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 
    6.4171e+06, 6.4172e+06, 6.4172e+06, 6.4172e+06, 6.4173e+06, 6.4173e+06, 
    6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4177e+06, 6.4177e+06, 
    6.4178e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 6.4179e+06, 6.418e+06, 
    6.418e+06, 6.418e+06, 6.4181e+06, 6.4181e+06, 6.4181e+06, 6.4182e+06, 
    6.4182e+06, 6.4182e+06, 6.4183e+06, 6.4183e+06, 6.4183e+06, 6.4184e+06, 
    6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4185e+06, 6.4186e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 
    6.4188e+06, 6.4189e+06, 6.4189e+06, 6.4189e+06, 6.419e+06, 6.419e+06, 
    6.419e+06, 6.4191e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4193e+06, 6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4194e+06, 
    6.4195e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 6.4196e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 
    6.4199e+06, 6.4199e+06, 6.42e+06, 6.42e+06, 6.42e+06, 6.4201e+06, 
    6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 6.4203e+06, 
    6.4203e+06, 6.4204e+06, 6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 
    6.4205e+06, 6.4206e+06, 6.4206e+06, 6.4206e+06, 6.4207e+06, 6.4207e+06, 
    6.4208e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.4209e+06, 6.4209e+06, 
    6.421e+06, 6.421e+06, 6.421e+06, 6.4211e+06, 6.4211e+06, 6.4212e+06, 
    6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4213e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 
    6.4216e+06, 6.4217e+06, 6.4217e+06, 6.4217e+06, 6.4218e+06, 6.4218e+06, 
    6.4218e+06, 6.4219e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.422e+06, 
    6.422e+06, 6.4221e+06, 6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4222e+06, 
    6.4223e+06, 6.4223e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 
    6.4227e+06, 6.4227e+06, 6.4228e+06, 6.4228e+06, 6.4228e+06, 6.4229e+06, 
    6.4229e+06, 6.423e+06, 6.423e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 
    6.4231e+06, 6.4232e+06, 6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4233e+06, 
    6.4234e+06, 6.4234e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 6.4236e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 
    6.4238e+06, 6.4238e+06, 6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 
    6.424e+06, 6.4241e+06, 6.4241e+06, 6.4241e+06, 6.4242e+06, 6.4242e+06, 
    6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4244e+06, 6.4244e+06, 
    6.4245e+06, 6.4245e+06, 6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4246e+06, 
    6.4247e+06, 6.4247e+06, 6.4248e+06, 6.4248e+06, 6.4248e+06, 6.4249e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 
    6.4251e+06, 6.4252e+06, 6.4252e+06, 6.4252e+06, 6.4253e+06, 6.4253e+06, 
    6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4256e+06, 6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4257e+06, 
    6.4258e+06, 6.4258e+06, 6.4259e+06, 6.4259e+06, 6.4259e+06, 6.426e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 
    6.4262e+06, 6.4263e+06, 6.4263e+06, 6.4263e+06, 6.4264e+06, 6.4264e+06, 
    6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 6.4266e+06, 6.4266e+06, 
    6.4267e+06, 6.4267e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4268e+06, 
    6.4269e+06, 6.4269e+06, 6.427e+06, 6.427e+06, 6.427e+06, 6.4271e+06, 
    6.4271e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4275e+06, 
    6.4275e+06, 6.4276e+06, 6.4276e+06, 6.4277e+06, 6.4277e+06, 6.4277e+06, 
    6.4278e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.428e+06, 6.4281e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 
    6.4282e+06, 6.4283e+06, 6.4283e+06, 6.4283e+06, 6.4284e+06, 6.4284e+06, 
    6.4284e+06, 6.4285e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4286e+06, 
    6.4287e+06, 6.4287e+06, 6.4287e+06, 6.4288e+06, 6.4288e+06, 6.4289e+06, 
    6.4289e+06, 6.4289e+06, 6.429e+06, 6.429e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 
    6.4293e+06, 6.4294e+06, 6.4294e+06, 6.4295e+06, 6.4295e+06, 6.4295e+06, 
    6.4296e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 6.4298e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.4299e+06, 6.4299e+06, 6.43e+06, 
    6.43e+06, 6.4301e+06, 6.4301e+06, 6.4301e+06, 6.4302e+06, 6.4302e+06, 
    6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4304e+06, 6.4305e+06, 6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4306e+06, 
    6.4307e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 6.4308e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 
    6.4311e+06, 6.4311e+06, 6.4312e+06, 6.4312e+06, 6.4313e+06, 6.4313e+06, 
    6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4317e+06, 
    6.4318e+06, 6.4318e+06, 6.4319e+06, 6.4319e+06, 6.4319e+06, 6.432e+06, 
    6.432e+06, 6.432e+06, 6.4321e+06, 6.4321e+06, 6.4322e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 
    6.4324e+06, 6.4325e+06, 6.4325e+06, 6.4326e+06, 6.4326e+06, 6.4326e+06, 
    6.4327e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.4329e+06, 6.433e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 
    6.4331e+06, 6.4331e+06, 6.4332e+06, 6.4332e+06, 6.4332e+06, 6.4333e+06, 
    6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4335e+06, 
    6.4335e+06, 6.4336e+06, 6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4337e+06, 
    6.4338e+06, 6.4338e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 6.434e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4342e+06, 
    6.4342e+06, 6.4343e+06, 6.4343e+06, 6.4343e+06, 6.4344e+06, 6.4344e+06, 
    6.4345e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 6.4346e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 
    6.4349e+06, 6.4349e+06, 6.435e+06, 6.435e+06, 6.435e+06, 6.4351e+06, 
    6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 6.4353e+06, 
    6.4353e+06, 6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4355e+06, 
    6.4356e+06, 6.4356e+06, 6.4356e+06, 6.4357e+06, 6.4357e+06, 6.4357e+06, 
    6.4358e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 
    6.436e+06, 6.436e+06, 6.4361e+06, 6.4361e+06, 6.4361e+06, 6.4362e+06, 
    6.4362e+06, 6.4363e+06, 6.4363e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4364e+06, 6.4365e+06, 6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4366e+06, 
    6.4367e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 6.4368e+06, 6.4368e+06, 
    6.4369e+06, 6.4369e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 
    6.4371e+06, 6.4371e+06, 6.4372e+06, 6.4372e+06, 6.4372e+06, 6.4373e+06, 
    6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 6.4375e+06, 6.4375e+06, 
    6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4377e+06, 
    6.4377e+06, 6.4378e+06, 6.4378e+06, 6.4379e+06, 6.4379e+06, 6.4379e+06, 
    6.438e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 6.4381e+06, 6.4382e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 
    6.4384e+06, 6.4385e+06, 6.4385e+06, 6.4385e+06, 6.4386e+06, 6.4386e+06, 
    6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.439e+06, 
    6.4391e+06, 6.4391e+06, 6.4392e+06, 6.4392e+06, 6.4392e+06, 6.4393e+06, 
    6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4394e+06, 6.4394e+06, 6.4395e+06, 
    6.4395e+06, 6.4396e+06, 6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4397e+06, 
    6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 6.4399e+06, 6.4399e+06, 
    6.44e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4401e+06, 
    6.4402e+06, 6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 
    6.4404e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 6.4406e+06, 6.4406e+06, 
    6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4408e+06, 
    6.4408e+06, 6.4409e+06, 6.4409e+06, 6.441e+06, 6.441e+06, 6.441e+06, 
    6.4411e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 6.4412e+06, 6.4413e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 
    6.4415e+06, 6.4416e+06, 6.4416e+06, 6.4416e+06, 6.4417e+06, 6.4417e+06, 
    6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.442e+06, 6.442e+06, 6.4421e+06, 6.4421e+06, 6.4421e+06, 
    6.4422e+06, 6.4422e+06, 6.4423e+06, 6.4423e+06, 6.4423e+06, 6.4424e+06, 
    6.4424e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4426e+06, 6.4427e+06, 6.4427e+06, 6.4427e+06, 6.4428e+06, 6.4428e+06, 
    6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 6.443e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4432e+06, 
    6.4433e+06, 6.4433e+06, 6.4434e+06, 6.4434e+06, 6.4434e+06, 6.4435e+06, 
    6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4437e+06, 6.4438e+06, 6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 
    6.4439e+06, 6.444e+06, 6.444e+06, 6.4441e+06, 6.4441e+06, 6.4441e+06, 
    6.4442e+06, 6.4442e+06, 6.4442e+06 ;

 bangle_L1 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle =
  0.016718, 0.016852, 0.017001, 0.017179, 0.01739, 0.017619, 0.017865, 
    0.018113, 0.018368, 0.018649, 0.018947, 0.019248, 0.019549, 0.019851, 
    0.020152, 0.020453, 0.020723, 0.020983, 0.021224, 0.02145, 0.021662, 
    0.021837, 0.021995, 0.0221, 0.022208, 0.022319, 0.022431, 0.022541, 
    0.022629, 0.022716, 0.022803, 0.022899, 0.022999, 0.023103, 0.023203, 
    0.023296, 0.023372, 0.023442, 0.023487, 0.023527, 0.023554, 0.023578, 
    0.0236, 0.023595, 0.023582, 0.023553, 0.023522, 0.023488, 0.023466, 
    0.023443, 0.02342, 0.023396, 0.023372, 0.023346, 0.023321, 0.023301, 
    0.023285, 0.023273, 0.023284, 0.0233, 0.023316, 0.02333, 0.023342, 
    0.023331, 0.023312, 0.023286, 0.023263, 0.023245, 0.023228, 0.023209, 
    0.02318, 0.023147, 0.023109, 0.02308, 0.023055, 0.023048, 0.023045, 
    0.023048, 0.02305, 0.02305, 0.023051, 0.02306, 0.023089, 0.023127, 
    0.023171, 0.023203, 0.023232, 0.023259, 0.023284, 0.023309, 0.023337, 
    0.023366, 0.023397, 0.023423, 0.023444, 0.023459, 0.023473, 0.023483, 
    0.023494, 0.023503, 0.023507, 0.02351, 0.023515, 0.023519, 0.023525, 
    0.023529, 0.023533, 0.023531, 0.023526, 0.023517, 0.023513, 0.023511, 
    0.02351, 0.023505, 0.023493, 0.023478, 0.023462, 0.023443, 0.023423, 
    0.023401, 0.02338, 0.023361, 0.023351, 0.023342, 0.023334, 0.023327, 
    0.023321, 0.023327, 0.023334, 0.023341, 0.023349, 0.023356, 0.02337, 
    0.023386, 0.023405, 0.023423, 0.023441, 0.02346, 0.023478, 0.023492, 
    0.023507, 0.023522, 0.02354, 0.023559, 0.023574, 0.023591, 0.023611, 
    0.023635, 0.02366, 0.023686, 0.02371, 0.02373, 0.023763, 0.023803, 
    0.023851, 0.023897, 0.023934, 0.023982, 0.024036, 0.024096, 0.024154, 
    0.024207, 0.024256, 0.024302, 0.024348, 0.024393, 0.024436, 0.024479, 
    0.024522, 0.024568, 0.024614, 0.024652, 0.024688, 0.024724, 0.024762, 
    0.024802, 0.024846, 0.024894, 0.024949, 0.025003, 0.025057, 0.025111, 
    0.025169, 0.025233, 0.025298, 0.025364, 0.025408, 0.025446, 0.025476, 
    0.025487, 0.025489, 0.025428, 0.02535, 0.025231, 0.025113, 0.024996, 
    0.024862, 0.024724, 0.024574, 0.024431, 0.024294, 0.024187, 0.024083, 
    0.023971, 0.023857, 0.023742, 0.023623, 0.023499, 0.023352, 0.023204, 
    0.023055, 0.022906, 0.022753, 0.022574, 0.022377, 0.022156, 0.021965, 
    0.021785, 0.021608, 0.021428, 0.021245, 0.021053, 0.020858, 0.020655, 
    0.020456, 0.020267, 0.020092, 0.019925, 0.019811, 0.019708, 0.019628, 
    0.019582, 0.019559, 0.019539, 0.019518, 0.019494, 0.019472, 0.019451, 
    0.019406, 0.019349, 0.019258, 0.01916, 0.019055, 0.01897, 0.018886, 
    0.018788, 0.018696, 0.018611, 0.018527, 0.018442, 0.01834, 0.018264, 
    0.018223, 0.018205, 0.018191, 0.018136, 0.01807, 0.017985, 0.017913, 
    0.017847, 0.017749, 0.017665, 0.017611, 0.017562, 0.017516, 0.017454, 
    0.017394, 0.01734, 0.017289, 0.017242, 0.017195, 0.01715, 0.017109, 
    0.01707, 0.017032, 0.016995, 0.016962, 0.016949, 0.016947, 0.016957, 
    0.016973, 0.016987, 0.016989, 0.017005, 0.017039, 0.017079, 0.017121, 
    0.017168, 0.017217, 0.017269, 0.017302, 0.017328, 0.017347, 0.017371, 
    0.017402, 0.017449, 0.017503, 0.017545, 0.0176, 0.017679, 0.017726, 
    0.017755, 0.017787, 0.017814, 0.017827, 0.017834, 0.017837, 0.017837, 
    0.017836, 0.017827, 0.017817, 0.017807, 0.017794, 0.017781, 0.017769, 
    0.017757, 0.017744, 0.017734, 0.017727, 0.017729, 0.017737, 0.017749, 
    0.017752, 0.017752, 0.017742, 0.017728, 0.017711, 0.017677, 0.017637, 
    0.017594, 0.017551, 0.01751, 0.017471, 0.017432, 0.017394, 0.017357, 
    0.017321, 0.01729, 0.017263, 0.017244, 0.017233, 0.017237, 0.017259, 
    0.017291, 0.017329, 0.017369, 0.01741, 0.017451, 0.017492, 0.017539, 
    0.017585, 0.017629, 0.017668, 0.017704, 0.017737, 0.017767, 0.017789, 
    0.017805, 0.017815, 0.017822, 0.017828, 0.017842, 0.017856, 0.017871, 
    0.017902, 0.01794, 0.017996, 0.01805, 0.018102, 0.01815, 0.018195, 
    0.018238, 0.018281, 0.018322, 0.01836, 0.018397, 0.018428, 0.018458, 
    0.018482, 0.018496, 0.018502, 0.018502, 0.018501, 0.0185, 0.018499, 
    0.018497, 0.018495, 0.018491, 0.018485, 0.018482, 0.018481, 0.018481, 
    0.018482, 0.018482, 0.018481, 0.018477, 0.018463, 0.018448, 0.018429, 
    0.018411, 0.018391, 0.018371, 0.018351, 0.018332, 0.018313, 0.018295, 
    0.018276, 0.018256, 0.018242, 0.018231, 0.018222, 0.018211, 0.018198, 
    0.018197, 0.018196, 0.018198, 0.018193, 0.018184, 0.018175, 0.018167, 
    0.018161, 0.018154, 0.018146, 0.018136, 0.018125, 0.018118, 0.018111, 
    0.018105, 0.018097, 0.018089, 0.018086, 0.018085, 0.018086, 0.018087, 
    0.018089, 0.018095, 0.018104, 0.018116, 0.018127, 0.018136, 0.018139, 
    0.018138, 0.018131, 0.018124, 0.018117, 0.018114, 0.018111, 0.018105, 
    0.018097, 0.018086, 0.018081, 0.018073, 0.018059, 0.018047, 0.018035, 
    0.018037, 0.018039, 0.018038, 0.018032, 0.018024, 0.018027, 0.018032, 
    0.018041, 0.018044, 0.018042, 0.018034, 0.018024, 0.018017, 0.018007, 
    0.017994, 0.017986, 0.017978, 0.017972, 0.017963, 0.017951, 0.017944, 
    0.017937, 0.017938, 0.017943, 0.017954, 0.017972, 0.017994, 0.018011, 
    0.018029, 0.018047, 0.018067, 0.018088, 0.018106, 0.018122, 0.018132, 
    0.018139, 0.018146, 0.018151, 0.018155, 0.018154, 0.018154, 0.018156, 
    0.018156, 0.018154, 0.018144, 0.018135, 0.018127, 0.018129, 0.018133, 
    0.018138, 0.018143, 0.018147, 0.018152, 0.018157, 0.018159, 0.018164, 
    0.018171, 0.018178, 0.018184, 0.018183, 0.01818, 0.018177, 0.018171, 
    0.018163, 0.018156, 0.018149, 0.018143, 0.018134, 0.018124, 0.018111, 
    0.018099, 0.018091, 0.018087, 0.018085, 0.018082, 0.018078, 0.018073, 
    0.018068, 0.018064, 0.01806, 0.018056, 0.018053, 0.018049, 0.018044, 
    0.018036, 0.018028, 0.018019, 0.018011, 0.018003, 0.017995, 0.017986, 
    0.017979, 0.017971, 0.017963, 0.017955, 0.017948, 0.017941, 0.017934, 
    0.017927, 0.017921, 0.017914, 0.017908, 0.017901, 0.017895, 0.017891, 
    0.017888, 0.017885, 0.017881, 0.017877, 0.017875, 0.017874, 0.017876, 
    0.017879, 0.017883, 0.017888, 0.017893, 0.017897, 0.017901, 0.017905, 
    0.017908, 0.017912, 0.017918, 0.017924, 0.01793, 0.017931, 0.017926, 
    0.01792, 0.017913, 0.017911, 0.017906, 0.017898, 0.017889, 0.01788, 
    0.01787, 0.01786, 0.01785, 0.017839, 0.017827, 0.017816, 0.017805, 
    0.017795, 0.017785, 0.017775, 0.017761, 0.017749, 0.017737, 0.017725, 
    0.017712, 0.017696, 0.017679, 0.01766, 0.017639, 0.017615, 0.017592, 
    0.017569, 0.017545, 0.017522, 0.0175, 0.01748, 0.017461, 0.017443, 
    0.017427, 0.017414, 0.017408, 0.017403, 0.017396, 0.017389, 0.017379, 
    0.017375, 0.017373, 0.017372, 0.017371, 0.01737, 0.017369, 0.017369, 
    0.017368, 0.017367, 0.017365, 0.017363, 0.01736, 0.017354, 0.017347, 
    0.017336, 0.017323, 0.01731, 0.017297, 0.017284, 0.017272, 0.01726, 
    0.01725, 0.017243, 0.017236, 0.017231, 0.017227, 0.017223, 0.017221, 
    0.017218, 0.017214, 0.01721, 0.017208, 0.017206, 0.017205, 0.017206, 
    0.017208, 0.017211, 0.017212, 0.017213, 0.017211, 0.017209, 0.017208, 
    0.017208, 0.017208, 0.017208, 0.017209, 0.017209, 0.017205, 0.017198, 
    0.01719, 0.017186, 0.017188, 0.017191, 0.017195, 0.017204, 0.017215, 
    0.017232, 0.017251, 0.01727, 0.017291, 0.017312, 0.017332, 0.017353, 
    0.017373, 0.017394, 0.017416, 0.017436, 0.017454, 0.01747, 0.017482, 
    0.017492, 0.017497, 0.017501, 0.017502, 0.017504, 0.017507, 0.017507, 
    0.017506, 0.017501, 0.017492, 0.017481, 0.017467, 0.017453, 0.017438, 
    0.017424, 0.017412, 0.017407, 0.017402, 0.017396, 0.017387, 0.017377, 
    0.01737, 0.017364, 0.017357, 0.017347, 0.017335, 0.017323, 0.017312, 
    0.017304, 0.017294, 0.017284, 0.017272, 0.017259, 0.017246, 0.017233, 
    0.017221, 0.017209, 0.017199, 0.017191, 0.017185, 0.01718, 0.017177, 
    0.017174, 0.017168, 0.017163, 0.01716, 0.017158, 0.017156, 0.017157, 
    0.017161, 0.017169, 0.017177, 0.017187, 0.017196, 0.017205, 0.017213, 
    0.017222, 0.017231, 0.017244, 0.017257, 0.01727, 0.017282, 0.017293, 
    0.017304, 0.017317, 0.017332, 0.017347, 0.017362, 0.017381, 0.017402, 
    0.017433, 0.017466, 0.017501, 0.017538, 0.017577, 0.017625, 0.017674, 
    0.017723, 0.017771, 0.017819, 0.017857, 0.017893, 0.017924, 0.017954, 
    0.017985, 0.018018, 0.018049, 0.018078, 0.018103, 0.018124, 0.018144, 
    0.018164, 0.018185, 0.018206, 0.018227, 0.018244, 0.01826, 0.018273, 
    0.018286, 0.018297, 0.018306, 0.018314, 0.01832, 0.018323, 0.018325, 
    0.018326, 0.018324, 0.018315, 0.018303, 0.018289, 0.018271, 0.01825, 
    0.018222, 0.01819, 0.018153, 0.018109, 0.018062, 0.018011, 0.017963, 
    0.017918, 0.017872, 0.017824, 0.017767, 0.01771, 0.017652, 0.017594, 
    0.017535, 0.017477, 0.017417, 0.017356, 0.017289, 0.017219, 0.017147, 
    0.017074, 0.016998, 0.016922, 0.016844, 0.016764, 0.016684, 0.016605, 
    0.016525, 0.016442, 0.016357, 0.016273, 0.016191, 0.016111, 0.016032, 
    0.015949, 0.015865, 0.015785, 0.015707, 0.015631, 0.015556, 0.015482, 
    0.015416, 0.015353, 0.015292, 0.015234, 0.015177, 0.015134, 0.015093, 
    0.01506, 0.015026, 0.014992, 0.01496, 0.014929, 0.014899, 0.01487, 
    0.014842, 0.014821, 0.014802, 0.014786, 0.014772, 0.01476, 0.014749, 
    0.01474, 0.014734, 0.014729, 0.014724, 0.014719, 0.014715, 0.014713, 
    0.01471, 0.014708, 0.014704, 0.0147, 0.014695, 0.014689, 0.014681, 
    0.014671, 0.014661, 0.014652, 0.014643, 0.014634, 0.014621, 0.014608, 
    0.014597, 0.014585, 0.014569, 0.014551, 0.014532, 0.014518, 0.014503, 
    0.014488, 0.014472, 0.014456, 0.014443, 0.014431, 0.01442, 0.014409, 
    0.014398, 0.014385, 0.014372, 0.014357, 0.014343, 0.014328, 0.014315, 
    0.014303, 0.01429, 0.014275, 0.014258, 0.014239, 0.01422, 0.014203, 
    0.014186, 0.014169, 0.014153, 0.014138, 0.014122, 0.014105, 0.014086, 
    0.01407, 0.014056, 0.014046, 0.014035, 0.014024, 0.014016, 0.014009, 
    0.014001, 0.013993, 0.013986, 0.013981, 0.013977, 0.013974, 0.01397, 
    0.013965, 0.013959, 0.013953, 0.013946, 0.01394, 0.013935, 0.01393, 
    0.013926, 0.013922, 0.013917, 0.013908, 0.013902, 0.013897, 0.013894, 
    0.013891, 0.013889, 0.013888, 0.013885, 0.013885, 0.013887, 0.013887, 
    0.013889, 0.013891, 0.013895, 0.013899, 0.013892, 0.013885, 0.013879, 
    0.013876, 0.013873, 0.013866, 0.013858, 0.013852, 0.013847, 0.013842, 
    0.013837, 0.013834, 0.013834, 0.013836, 0.013838, 0.01384, 0.013842, 
    0.013843, 0.013845, 0.013849, 0.013852, 0.013855, 0.013858, 0.013861, 
    0.013864, 0.013865, 0.013866, 0.013866, 0.013867, 0.013869, 0.013871, 
    0.013873, 0.013874, 0.013874, 0.013875, 0.013875, 0.013875, 0.013876, 
    0.013879, 0.013886, 0.013891, 0.013895, 0.013896, 0.013899, 0.013905, 
    0.013909, 0.01391, 0.013913, 0.013915, 0.013917, 0.013917, 0.013914, 
    0.01391, 0.013906, 0.013902, 0.013899, 0.013896, 0.013892, 0.013886, 
    0.013876, 0.013865, 0.013853, 0.013842, 0.013831, 0.01382, 0.01381, 
    0.0138, 0.013789, 0.013778, 0.013765, 0.013754, 0.013744, 0.013736, 
    0.013729, 0.013719, 0.013711, 0.013704, 0.013695, 0.013686, 0.013679, 
    0.013672, 0.013664, 0.013655, 0.013647, 0.013637, 0.013626, 0.013616, 
    0.013606, 0.013594, 0.013582, 0.01357, 0.013559, 0.013547, 0.013535, 
    0.013524, 0.013513, 0.013502, 0.013495, 0.013491, 0.013487, 0.013482, 
    0.013483, 0.013482, 0.013479, 0.01348, 0.013481, 0.013483, 0.013484, 
    0.013481, 0.013477, 0.013471, 0.013466, 0.013461, 0.013459, 0.013455, 
    0.01345, 0.013447, 0.013443, 0.013438, 0.013432, 0.013427, 0.013424, 
    0.013423, 0.013428, 0.013429, 0.013429, 0.013428, 0.013427, 0.013428, 
    0.013429, 0.013429, 0.013429, 0.013429, 0.01343, 0.013431, 0.013432, 
    0.01343, 0.013428, 0.01343, 0.01343, 0.013429, 0.013431, 0.013434, 
    0.013427, 0.013422, 0.013418, 0.013418, 0.013418, 0.013417, 0.013415, 
    0.013411, 0.013405, 0.013397, 0.01339, 0.013383, 0.013374, 0.013367, 
    0.01336, 0.013355, 0.013348, 0.013339, 0.013329, 0.013317, 0.013308, 
    0.013299, 0.013289, 0.013277, 0.013266, 0.013256, 0.013246, 0.013237, 
    0.013227, 0.013217, 0.013205, 0.013193, 0.013183, 0.013171, 0.013157, 
    0.013144, 0.01313, 0.013114, 0.013101, 0.013092, 0.013081, 0.013068, 
    0.013057, 0.013046, 0.013036, 0.013028, 0.013022, 0.013017, 0.013013, 
    0.01301, 0.013007, 0.013005, 0.013, 0.012995, 0.01299, 0.012985, 0.01298, 
    0.012975, 0.012971, 0.012966, 0.012964, 0.012962, 0.01296, 0.012957, 
    0.012956, 0.012954, 0.012951, 0.012949, 0.012947, 0.012947, 0.012949, 
    0.012951, 0.012952, 0.012952, 0.012953, 0.012955, 0.012956, 0.012957, 
    0.012958, 0.012961, 0.012963, 0.012967, 0.012971, 0.012977, 0.012977, 
    0.012977, 0.012978, 0.012977, 0.012973, 0.012969, 0.012964, 0.01296, 
    0.012957, 0.012955, 0.012952, 0.012949, 0.012945, 0.012941, 0.012936, 
    0.012931, 0.012927, 0.012924, 0.012921, 0.012918, 0.012916, 0.012913, 
    0.012908, 0.012904, 0.0129, 0.012896, 0.012893, 0.012888, 0.012884, 
    0.012882, 0.01288, 0.012878, 0.012875, 0.012872, 0.012866, 0.012857, 
    0.012846, 0.012837, 0.012829, 0.012823, 0.012814, 0.012805, 0.012794, 
    0.012785, 0.012778, 0.01277, 0.012763, 0.012753, 0.012744, 0.012739, 
    0.012734, 0.01273, 0.012726, 0.012722, 0.012718, 0.012712, 0.012705, 
    0.012697, 0.012689, 0.012683, 0.012679, 0.012676, 0.01267, 0.012663, 
    0.012657, 0.012651, 0.012646, 0.012639, 0.012631, 0.012623, 0.012615, 
    0.012607, 0.012602, 0.012599, 0.012597, 0.012596, 0.012596, 0.012595, 
    0.012594, 0.012597, 0.012601, 0.012607, 0.012612, 0.012617, 0.012621, 
    0.012625, 0.012628, 0.01263, 0.012631, 0.012633, 0.012634, 0.012635, 
    0.012636, 0.012638, 0.01264, 0.012643, 0.012645, 0.012648, 0.012651, 
    0.012652, 0.012652, 0.01265, 0.012648, 0.012646, 0.012644, 0.012642, 
    0.012639, 0.012636, 0.012633, 0.012629, 0.012625, 0.01262, 0.012616, 
    0.012611, 0.012607, 0.012602, 0.012596, 0.01259, 0.012584, 0.012579, 
    0.012573, 0.012569, 0.012564, 0.01256, 0.012555, 0.012551, 0.012546, 
    0.01254, 0.012534, 0.012527, 0.012519, 0.012511, 0.012503, 0.012496, 
    0.012487, 0.012477, 0.012467, 0.012457, 0.012452, 0.012447, 0.012443, 
    0.01244, 0.012437, 0.012435, 0.012432, 0.012428, 0.012424, 0.012419, 
    0.012415, 0.012411, 0.012406, 0.012399, 0.012391, 0.012381, 0.012373, 
    0.012366, 0.01236, 0.012355, 0.012348, 0.012341, 0.012335, 0.01233, 
    0.012325, 0.01232, 0.012314, 0.012309, 0.012306, 0.012304, 0.0123, 
    0.012295, 0.01229, 0.012286, 0.012283, 0.012279, 0.012275, 0.012273, 
    0.012271, 0.012269, 0.012267, 0.012264, 0.012256, 0.012249, 0.012245, 
    0.012241, 0.012237, 0.012232, 0.012226, 0.012218, 0.012211, 0.012206, 
    0.012204, 0.012203, 0.012203, 0.012201, 0.012198, 0.012191, 0.012185, 
    0.012181, 0.012176, 0.01217, 0.012165, 0.012159, 0.012153, 0.012147, 
    0.012139, 0.012131, 0.012124, 0.012119, 0.012114, 0.012108, 0.012101, 
    0.012093, 0.012088, 0.012081, 0.012071, 0.012058, 0.012043, 0.012031, 
    0.01202, 0.01201, 0.012, 0.011988, 0.011977, 0.011967, 0.011959, 
    0.011951, 0.011942, 0.011934, 0.011925, 0.011917, 0.011908, 0.011898, 
    0.011888, 0.011878, 0.011868, 0.011859, 0.01185, 0.01184, 0.01183, 
    0.011821, 0.011813, 0.011806, 0.011799, 0.011792, 0.011784, 0.011778, 
    0.011773, 0.011768, 0.011764, 0.01176, 0.011755, 0.01175, 0.011747, 
    0.011746, 0.011745, 0.011745, 0.011744, 0.011743, 0.01174, 0.011738, 
    0.011736, 0.011735, 0.011735, 0.011735, 0.011734, 0.011733, 0.01173, 
    0.011726, 0.011723, 0.011721, 0.011721, 0.011723, 0.011723, 0.011721, 
    0.01172, 0.011719, 0.011717, 0.011715, 0.011714, 0.011711, 0.011708, 
    0.011707, 0.011706, 0.011705, 0.011702, 0.011698, 0.011694, 0.011691, 
    0.011687, 0.011681, 0.011675, 0.01167, 0.011666, 0.011663, 0.011658, 
    0.011652, 0.011647, 0.011642, 0.011639, 0.011636, 0.011633, 0.011629, 
    0.011625, 0.011622, 0.011619, 0.011616, 0.01161, 0.011605, 0.011602, 
    0.011598, 0.011592, 0.011589, 0.011586, 0.011581, 0.011577, 0.011574, 
    0.011572, 0.01157, 0.011569, 0.011567, 0.011565, 0.011564, 0.011563, 
    0.01156, 0.011558, 0.011556, 0.011554, 0.011554, 0.011553, 0.011552, 
    0.011551, 0.011549, 0.011546, 0.011544, 0.011542, 0.01154, 0.011538, 
    0.011535, 0.011529, 0.011524, 0.011519, 0.011514, 0.01151, 0.011506, 
    0.011501, 0.011497, 0.011492, 0.011486, 0.011478, 0.011471, 0.011465, 
    0.01146, 0.011457, 0.011451, 0.011445, 0.011438, 0.011431, 0.011424, 
    0.011415, 0.011406, 0.011397, 0.01139, 0.011385, 0.01138, 0.011376, 
    0.011371, 0.011365, 0.01136, 0.011356, 0.011351, 0.011348, 0.011345, 
    0.011344, 0.011341, 0.011338, 0.011335, 0.011332, 0.011328, 0.011324, 
    0.011319, 0.011314, 0.011309, 0.011303, 0.011297, 0.011292, 0.011289, 
    0.011286, 0.011285, 0.011283, 0.011281, 0.011276, 0.011272, 0.011269, 
    0.011267, 0.011266, 0.011267, 0.011268, 0.011268, 0.011267, 0.011265, 
    0.011262, 0.011258, 0.011254, 0.011251, 0.011247, 0.011244, 0.01124, 
    0.011237, 0.011233, 0.011228, 0.011224, 0.011219, 0.011215, 0.011211, 
    0.011208, 0.011205, 0.011203, 0.011204, 0.011204, 0.011204, 0.011203, 
    0.011202, 0.011199, 0.011195, 0.011194, 0.011192, 0.011192, 0.011191, 
    0.01119, 0.011189, 0.011187, 0.011184, 0.011181, 0.011178, 0.011174, 
    0.011171, 0.011169, 0.011167, 0.011165, 0.011161, 0.011158, 0.011154, 
    0.011151, 0.011148, 0.011142, 0.011137, 0.011135, 0.011135, 0.011135, 
    0.011135, 0.011134, 0.011133, 0.011132, 0.011131, 0.011129, 0.011127, 
    0.011125, 0.011123, 0.011122, 0.011124, 0.011125, 0.011127, 0.011128, 
    0.011126, 0.011124, 0.011121, 0.01112, 0.011121, 0.011122, 0.011122, 
    0.011121, 0.011119, 0.011117, 0.011113, 0.01111, 0.011108, 0.011105, 
    0.011103, 0.011101, 0.011098, 0.011095, 0.01109, 0.011086, 0.011082, 
    0.011075, 0.011067, 0.011061, 0.011055, 0.011051, 0.011047, 0.011043, 
    0.01104, 0.011037, 0.011032, 0.011027, 0.01102, 0.011016, 0.011012, 
    0.011008, 0.011002, 0.010995, 0.010989, 0.010982, 0.010976, 0.010968, 
    0.01096, 0.010951, 0.010942, 0.010934, 0.010926, 0.010918, 0.010911, 
    0.010903, 0.010895, 0.010888, 0.010881, 0.010875, 0.01087, 0.010864, 
    0.010858, 0.010854, 0.010851, 0.010849, 0.010845, 0.010842, 0.010837, 
    0.010831, 0.010824, 0.010819, 0.010812, 0.010804, 0.010798, 0.010794, 
    0.010788, 0.010783, 0.010775, 0.010768, 0.010761, 0.010756, 0.010752, 
    0.010748, 0.010745, 0.010741, 0.01074, 0.010739, 0.010737, 0.010736, 
    0.010735, 0.010734, 0.010734, 0.010735, 0.010737, 0.010738, 0.010737, 
    0.010735, 0.010731, 0.010727, 0.010725, 0.010722, 0.010721, 0.010719, 
    0.010716, 0.010709, 0.010702, 0.010696, 0.010692, 0.01069, 0.010692, 
    0.010695, 0.010697, 0.010696, 0.010694, 0.010693, 0.010691, 0.010689, 
    0.01069, 0.010691, 0.010691, 0.010691, 0.01069, 0.010687, 0.010684, 
    0.01068, 0.010676, 0.010673, 0.01067, 0.010668, 0.010663, 0.010658, 
    0.010653, 0.010647, 0.010642, 0.010641, 0.01064, 0.010641, 0.010641, 
    0.010641, 0.010637, 0.010633, 0.010631, 0.010631, 0.010632, 0.010634, 
    0.010635, 0.010633, 0.010628, 0.010618, 0.010612, 0.010607, 0.010603, 
    0.0106, 0.010599, 0.010596, 0.010591, 0.010587, 0.010582, 0.010577, 
    0.010572, 0.010567, 0.010563, 0.010558, 0.010553, 0.010547, 0.010542, 
    0.010536, 0.01053, 0.010524, 0.010518, 0.010512, 0.010505, 0.010497, 
    0.010488, 0.010479, 0.01047, 0.010464, 0.010458, 0.010452, 0.010446, 
    0.010439, 0.010431, 0.010423, 0.010412, 0.010402, 0.010394, 0.010387, 
    0.01038, 0.010369, 0.010358, 0.010345, 0.010333, 0.010321, 0.010311, 
    0.010301, 0.010292, 0.010283, 0.010274, 0.010266, 0.010259, 0.010252, 
    0.010245, 0.010238, 0.010231, 0.010224, 0.010218, 0.01021, 0.010202, 
    0.010196, 0.010189, 0.010183, 0.010178, 0.010174, 0.010169, 0.010162, 
    0.010156, 0.010148, 0.010141, 0.010134, 0.010128, 0.010124, 0.01012, 
    0.010115, 0.010111, 0.010108, 0.010103, 0.010102, 0.010103, 0.010105, 
    0.010107, 0.01011, 0.010112, 0.010112, 0.010113, 0.010113, 0.010114, 
    0.010114, 0.010115, 0.010117, 0.010119, 0.01012, 0.010121, 0.010122, 
    0.010123, 0.010123, 0.010124, 0.010126, 0.010128, 0.010129, 0.010131, 
    0.010132, 0.010132, 0.010134, 0.010136, 0.010139, 0.010142, 0.010146, 
    0.010149, 0.010151, 0.010154, 0.010156, 0.010158, 0.010159, 0.01016, 
    0.010163, 0.010163, 0.010162, 0.010159, 0.010156, 0.010153, 0.010152, 
    0.010152, 0.010152, 0.010151, 0.01015, 0.010149, 0.010148, 0.010147, 
    0.010146, 0.010145, 0.010144, 0.010143, 0.010144, 0.010144, 0.010143, 
    0.010143, 0.010143, 0.010142, 0.010142, 0.010143, 0.010143, 0.010141, 
    0.01014, 0.010138, 0.010135, 0.010133, 0.010131, 0.010129, 0.010126, 
    0.010123, 0.01012, 0.010115, 0.01011, 0.010106, 0.010105, 0.010104, 
    0.010105, 0.010106, 0.010106, 0.010103, 0.010099, 0.010097, 0.010095, 
    0.010093, 0.010092, 0.010089, 0.010086, 0.010079, 0.010072, 0.010065, 
    0.010058, 0.010052, 0.010048, 0.010045, 0.010042, 0.010039, 0.010035, 
    0.010031, 0.010026, 0.010021, 0.010016, 0.010013, 0.010012, 0.010011, 
    0.010006, 0.01, 0.0099963, 0.0099919, 0.0099869, 0.0099846, 0.0099827, 
    0.0099798, 0.0099758, 0.0099705, 0.0099629, 0.0099545, 0.0099459, 
    0.0099387, 0.0099337, 0.0099277, 0.0099214, 0.0099155, 0.0099089, 
    0.0099006, 0.009894, 0.0098882, 0.0098872, 0.0098861, 0.0098846, 
    0.0098834, 0.0098824, 0.0098783, 0.0098739, 0.0098688, 0.0098633, 
    0.0098574, 0.0098547, 0.0098527, 0.0098521, 0.009849, 0.0098436, 
    0.009837, 0.0098304, 0.0098248, 0.0098198, 0.0098153, 0.0098113, 
    0.0098076, 0.0098038, 0.0097988, 0.0097921, 0.0097864, 0.0097813, 
    0.00978, 0.0097788, 0.0097776, 0.0097766, 0.0097756, 0.0097727, 
    0.0097701, 0.0097679, 0.0097669, 0.0097665, 0.0097674, 0.0097675, 
    0.0097657, 0.009763, 0.0097598, 0.0097534, 0.0097467, 0.0097396, 
    0.0097363, 0.009736, 0.0097321, 0.009727, 0.0097189, 0.0097102, 
    0.0097011, 0.0096947, 0.0096893, 0.0096859, 0.0096822, 0.0096781, 
    0.0096742, 0.00967, 0.0096644, 0.009659, 0.0096539, 0.0096525, 0.0096521, 
    0.0096508, 0.0096488, 0.0096458, 0.00964, 0.0096332, 0.0096273, 
    0.0096211, 0.0096144, 0.0096076, 0.0096007, 0.0095942, 0.0095878, 
    0.0095816, 0.0095759, 0.0095706, 0.0095653, 0.0095602, 0.009556, 
    0.0095524, 0.0095493, 0.0095417, 0.0095347, 0.0095329, 0.0095306, 
    0.0095278, 0.0095246, 0.0095215, 0.0095184, 0.0095154, 0.0095127, 
    0.0095107, 0.0095088, 0.0095059, 0.0095033, 0.0095012, 0.0094965, 
    0.0094908, 0.009484, 0.0094772, 0.0094703, 0.0094656, 0.009462, 
    0.0094606, 0.0094592, 0.0094578, 0.0094574, 0.0094576, 0.009456, 
    0.0094541, 0.0094516, 0.0094481, 0.0094441, 0.0094404, 0.0094366, 
    0.0094325, 0.009429, 0.0094259, 0.0094219, 0.0094175, 0.0094123, 
    0.0094079, 0.0094042, 0.0094017, 0.0093994, 0.0093972, 0.0093944, 
    0.0093909, 0.0093874, 0.0093841, 0.0093815, 0.0093799, 0.0093796, 
    0.0093789, 0.0093782, 0.0093791, 0.0093801, 0.0093815, 0.0093819, 
    0.0093819, 0.0093812, 0.0093799, 0.0093775, 0.0093739, 0.0093698, 
    0.0093656, 0.0093615, 0.0093578, 0.0093527, 0.0093467, 0.0093403, 
    0.0093343, 0.0093298, 0.0093257, 0.0093221, 0.0093185, 0.009315, 
    0.0093123, 0.0093093, 0.0093062, 0.0093021, 0.0092979, 0.0092943, 
    0.0092905, 0.0092864, 0.0092833, 0.0092804, 0.0092772, 0.0092734, 
    0.0092686, 0.009264, 0.0092596, 0.0092562, 0.0092524, 0.0092477, 
    0.0092427, 0.0092376, 0.0092324, 0.0092273, 0.0092222, 0.0092162, 
    0.0092097, 0.0092028, 0.0091952, 0.0091862, 0.0091781, 0.0091705, 
    0.009168, 0.0091661, 0.0091646, 0.0091628, 0.0091607, 0.0091575, 
    0.0091538, 0.0091491, 0.0091446, 0.0091405, 0.0091362, 0.0091322, 
    0.0091301, 0.0091275, 0.0091243, 0.0091215, 0.0091186, 0.0091145, 
    0.0091105, 0.0091067, 0.0091025, 0.0090982, 0.0090927, 0.0090876, 
    0.009083, 0.0090776, 0.0090719, 0.0090657, 0.0090595, 0.0090533, 
    0.0090474, 0.0090417, 0.0090383, 0.0090359, 0.0090353, 0.0090354, 
    0.009036, 0.009035, 0.0090335, 0.0090304, 0.0090273, 0.0090242, 
    0.0090207, 0.0090176, 0.0090159, 0.009014, 0.0090118, 0.009008, 
    0.0090035, 0.0089968, 0.0089898, 0.0089826, 0.0089771, 0.0089723, 
    0.0089701, 0.0089678, 0.0089655, 0.0089606, 0.008955, 0.0089515, 
    0.0089486, 0.0089468, 0.0089483, 0.0089512, 0.0089507, 0.00895, 
    0.0089493, 0.008948, 0.0089463, 0.0089453, 0.0089443, 0.008943, 
    0.0089415, 0.0089397, 0.0089388, 0.008938, 0.0089369, 0.0089359, 
    0.0089349, 0.0089331, 0.0089313, 0.0089297, 0.0089276, 0.0089249, 
    0.0089239, 0.0089235, 0.0089245, 0.0089262, 0.0089284, 0.0089305, 
    0.0089322, 0.0089315, 0.0089296, 0.0089261, 0.0089227, 0.0089196, 
    0.0089212, 0.00892, 0.0089147, 0.0089075, 0.0088994, 0.0088896, 
    0.0088812, 0.0088753, 0.0088701, 0.0088652, 0.008862, 0.0088585, 
    0.0088538, 0.0088487, 0.0088435, 0.008841, 0.0088388, 0.0088368, 
    0.008834, 0.0088305, 0.0088254, 0.00882, 0.0088145, 0.0088093, 0.0088044, 
    0.0088017, 0.0087993, 0.0087953, 0.0087915, 0.008788, 0.008784, 
    0.0087798, 0.0087752, 0.0087709, 0.0087671, 0.0087646, 0.0087623, 
    0.008759, 0.0087557, 0.0087525, 0.0087506, 0.0087492, 0.0087492, 
    0.0087489, 0.0087482, 0.008748, 0.0087482, 0.0087483, 0.008749, 
    0.0087514, 0.0087545, 0.0087581, 0.00876, 0.0087614, 0.008762, 0.0087614, 
    0.0087599, 0.00876, 0.0087606, 0.0087623, 0.0087629, 0.0087627, 
    0.0087614, 0.0087597, 0.0087564, 0.0087541, 0.0087527, 0.0087512, 
    0.0087498, 0.0087488, 0.0087482, 0.008748, 0.0087465, 0.0087445, 
    0.0087428, 0.0087411, 0.0087394, 0.0087385, 0.0087379, 0.0087375, 
    0.0087365, 0.0087342, 0.0087329, 0.008732, 0.0087308, 0.0087291, 
    0.0087264, 0.0087227, 0.0087186, 0.0087137, 0.0087088, 0.0087038, 
    0.0086995, 0.0086958, 0.0086928, 0.0086897, 0.0086852, 0.0086804, 
    0.0086754, 0.0086703, 0.0086653, 0.0086603, 0.0086552, 0.0086499, 
    0.0086442, 0.0086383, 0.0086323, 0.0086263, 0.0086202, 0.0086146, 
    0.0086095, 0.0086069, 0.0086043, 0.0086018, 0.008599, 0.008596, 0.008594, 
    0.0085923, 0.0085913, 0.0085892, 0.0085865, 0.0085819, 0.0085774, 
    0.0085735, 0.0085688, 0.0085636, 0.0085606, 0.0085581, 0.0085568, 
    0.0085554, 0.0085541, 0.0085489, 0.0085432, 0.008537, 0.0085318, 
    0.0085275, 0.0085236, 0.0085201, 0.0085182, 0.0085166, 0.0085154, 
    0.0085143, 0.0085133, 0.0085132, 0.0085132, 0.0085134, 0.0085125, 
    0.0085111, 0.0085086, 0.0085051, 0.0084998, 0.0084966, 0.0084942, 
    0.008491, 0.0084868, 0.0084808, 0.0084757, 0.0084711, 0.0084705, 
    0.0084707, 0.0084727, 0.0084734, 0.0084733, 0.0084743, 0.0084745, 
    0.0084724, 0.0084699, 0.008467, 0.0084647, 0.0084627, 0.0084621, 
    0.0084621, 0.0084626, 0.0084638, 0.0084653, 0.0084672, 0.008469, 
    0.0084707, 0.0084715, 0.0084719, 0.0084719, 0.0084709, 0.0084685, 
    0.0084671, 0.008466, 0.0084638, 0.0084611, 0.0084576, 0.0084536, 
    0.0084495, 0.0084462, 0.0084433, 0.0084412, 0.0084401, 0.0084394, 
    0.0084389, 0.0084376, 0.0084342, 0.0084308, 0.0084275, 0.0084242, 
    0.0084209, 0.0084179, 0.0084148, 0.0084117, 0.0084089, 0.0084058, 
    0.0084014, 0.0083974, 0.0083939, 0.0083888, 0.0083832, 0.0083766, 
    0.0083695, 0.0083619, 0.0083545, 0.0083472, 0.0083403, 0.0083339, 
    0.0083282, 0.0083232, 0.0083184, 0.0083128, 0.0083083, 0.0083054, 
    0.0083041, 0.0083034, 0.0083021, 0.0082999, 0.0082963, 0.0082925, 
    0.0082887, 0.0082838, 0.008278, 0.0082701, 0.008262, 0.0082538, 
    0.0082455, 0.0082372, 0.0082291, 0.0082211, 0.0082132, 0.0082052, 
    0.008197, 0.0081882, 0.0081811, 0.0081755, 0.008171, 0.0081671, 
    0.0081656, 0.0081636, 0.0081612, 0.0081591, 0.008157, 0.0081552, 
    0.0081535, 0.0081518, 0.0081499, 0.0081479, 0.0081446, 0.0081413, 
    0.008138, 0.0081335, 0.0081285, 0.0081234, 0.0081185, 0.0081137, 
    0.0081092, 0.0081049, 0.0081019, 0.0080992, 0.0080974, 0.008097, 
    0.0080975, 0.0080982, 0.008099, 0.0081001, 0.0081006, 0.0081006, 
    0.0080987, 0.0080969, 0.0080962, 0.0080955, 0.0080949, 0.0080926, 
    0.0080898, 0.0080861, 0.0080816, 0.0080762, 0.0080717, 0.0080675, 
    0.0080646, 0.0080624, 0.0080609, 0.0080595, 0.008058, 0.008057, 
    0.0080563, 0.0080561, 0.0080562, 0.0080564, 0.0080572, 0.0080572, 
    0.0080559, 0.0080557, 0.008056, 0.0080547, 0.0080532, 0.0080513, 
    0.0080495, 0.008048, 0.0080476, 0.0080471, 0.0080462, 0.0080455, 
    0.0080449, 0.0080454, 0.0080461, 0.008047, 0.0080478, 0.0080484, 
    0.0080478, 0.008047, 0.0080462, 0.0080449, 0.0080432, 0.0080427, 
    0.0080428, 0.0080445, 0.0080459, 0.0080468, 0.0080471, 0.008047, 
    0.0080456, 0.0080447, 0.0080444, 0.0080435, 0.0080424, 0.0080414, 
    0.0080397, 0.0080368, 0.0080344, 0.0080321, 0.0080312, 0.0080311, 
    0.0080328, 0.0080334, 0.0080334, 0.0080321, 0.0080304, 0.008028, 
    0.0080259, 0.0080239, 0.0080217, 0.0080193, 0.0080168, 0.0080142, 
    0.0080116, 0.008009, 0.0080069, 0.0080075, 0.0080084, 0.0080096, 
    0.0080107, 0.0080117, 0.0080125, 0.0080123, 0.008011, 0.00801, 0.008009, 
    0.0080071, 0.0080048, 0.0080021, 0.0079993, 0.0079967, 0.007994, 
    0.0079916, 0.0079895, 0.0079886, 0.0079883, 0.0079867, 0.0079844, 
    0.0079805, 0.0079759, 0.0079708, 0.0079666, 0.0079625, 0.007958, 
    0.0079536, 0.0079491, 0.0079443, 0.0079397, 0.0079357, 0.0079325, 
    0.0079301, 0.0079275, 0.0079248, 0.0079214, 0.0079177, 0.0079138, 
    0.0079102, 0.007907, 0.0079059, 0.0079045, 0.0079026, 0.0078997, 
    0.0078964, 0.0078918, 0.007888, 0.0078857, 0.0078845, 0.0078836, 
    0.0078815, 0.0078798, 0.0078787, 0.0078774, 0.0078761, 0.0078742, 
    0.0078724, 0.0078708, 0.0078692, 0.0078676, 0.0078669, 0.0078662, 
    0.0078653, 0.0078644, 0.0078634, 0.0078618, 0.0078604, 0.0078596, 
    0.0078586, 0.0078574, 0.0078556, 0.0078536, 0.0078509, 0.0078478, 
    0.0078444, 0.0078417, 0.0078392, 0.007837, 0.0078341, 0.0078303, 
    0.0078269, 0.0078238, 0.0078209, 0.0078182, 0.0078156, 0.0078132, 
    0.007811, 0.0078086, 0.0078063, 0.0078043, 0.0078021, 0.0077996, 
    0.0077968, 0.0077942, 0.0077923, 0.0077904, 0.0077885, 0.0077868, 
    0.0077846, 0.007781, 0.0077777, 0.0077747, 0.0077721, 0.0077693, 
    0.0077659, 0.0077625, 0.0077592, 0.0077561, 0.0077533, 0.0077514, 
    0.0077498, 0.0077487, 0.0077475, 0.0077459, 0.007742, 0.0077379, 
    0.0077337, 0.0077305, 0.0077275, 0.0077234, 0.007719, 0.0077139, 
    0.0077086, 0.0077032, 0.0076974, 0.0076916, 0.0076858, 0.0076793, 
    0.0076725, 0.007667, 0.0076617, 0.0076567, 0.0076522, 0.007648, 
    0.0076442, 0.0076408, 0.0076381, 0.0076363, 0.0076352, 0.007635, 
    0.0076349, 0.0076349, 0.0076341, 0.0076327, 0.0076297, 0.0076263, 
    0.0076218, 0.0076177, 0.0076141, 0.0076108, 0.0076075, 0.0076031, 
    0.007599, 0.0075951, 0.0075903, 0.0075853, 0.007581, 0.0075777, 
    0.0075758, 0.007574, 0.0075722, 0.0075704, 0.0075683, 0.007566, 
    0.0075645, 0.0075633, 0.0075631, 0.007563, 0.0075631, 0.0075628, 
    0.0075623, 0.0075602, 0.0075579, 0.007555, 0.0075518, 0.0075483, 
    0.0075454, 0.007542, 0.007537, 0.0075322, 0.0075275, 0.0075253, 
    0.0075239, 0.0075234, 0.0075232, 0.0075233, 0.007522, 0.0075205, 
    0.0075195, 0.0075182, 0.0075165, 0.0075169, 0.0075177, 0.0075152, 
    0.0075123, 0.0075087, 0.0075065, 0.0075049, 0.0075025, 0.0075008, 
    0.0075001, 0.0075011, 0.0075029, 0.0075045, 0.0075055, 0.0075052, 
    0.0075046, 0.0075038, 0.0075022, 0.0075006, 0.0074994, 0.0074981, 
    0.0074967, 0.0074942, 0.0074912, 0.0074865, 0.0074831, 0.0074809, 
    0.0074797, 0.0074784, 0.0074758, 0.0074732, 0.0074704, 0.0074679, 
    0.0074655, 0.007464, 0.0074626, 0.0074615, 0.0074614, 0.0074615, 
    0.0074607, 0.0074609, 0.0074624, 0.0074637, 0.0074648, 0.0074635, 
    0.0074629, 0.0074635, 0.0074618, 0.0074589, 0.0074538, 0.0074486, 
    0.0074434, 0.0074382, 0.0074329, 0.0074286, 0.0074247, 0.0074217, 
    0.0074187, 0.0074158, 0.0074134, 0.0074111, 0.0074092, 0.0074076, 
    0.0074062, 0.0074042, 0.0074017, 0.0073982, 0.0073964, 0.0073965, 
    0.0073979, 0.0073994, 0.0073987, 0.0073966, 0.0073927, 0.0073896, 
    0.0073869, 0.0073843, 0.0073821, 0.0073806, 0.0073788, 0.007377, 
    0.007374, 0.0073713, 0.0073692, 0.0073676, 0.0073662, 0.007366, 
    0.0073657, 0.0073648, 0.0073639, 0.0073631, 0.0073633, 0.0073637, 
    0.007364, 0.0073648, 0.0073659, 0.0073663, 0.0073664, 0.0073653, 
    0.0073641, 0.0073626, 0.0073615, 0.0073604, 0.0073596, 0.0073589, 
    0.0073582, 0.0073542, 0.0073493, 0.0073438, 0.0073396, 0.0073371, 
    0.0073361, 0.0073356, 0.0073352, 0.0073344, 0.0073327, 0.0073299, 
    0.0073266, 0.0073225, 0.0073188, 0.0073159, 0.0073127, 0.0073092, 
    0.0073051, 0.0073012, 0.0072982, 0.0072954, 0.0072929, 0.0072914, 
    0.0072898, 0.007288, 0.0072862, 0.0072845, 0.0072828, 0.0072815, 
    0.0072818, 0.0072824, 0.0072831, 0.0072835, 0.0072838, 0.0072838, 
    0.0072839, 0.007284, 0.007284, 0.0072841, 0.0072846, 0.0072853, 0.007286, 
    0.0072867, 0.0072873, 0.0072883, 0.0072898, 0.0072918, 0.0072942, 
    0.0072969, 0.0073012, 0.0073057, 0.0073108, 0.0073156, 0.0073204, 
    0.0073248, 0.0073286, 0.007331, 0.0073326, 0.0073337, 0.0073345, 
    0.0073352, 0.0073357, 0.0073364, 0.0073372, 0.0073393, 0.0073412, 
    0.0073422, 0.0073428, 0.0073431, 0.0073451, 0.0073474, 0.0073498, 
    0.0073522, 0.0073546, 0.007357, 0.0073594, 0.007362, 0.0073642, 
    0.0073657, 0.0073677, 0.0073698, 0.0073714, 0.0073729, 0.0073743, 
    0.0073753, 0.0073761, 0.007376, 0.0073752, 0.0073733, 0.0073712, 
    0.0073691, 0.0073679, 0.0073669, 0.0073663, 0.0073671, 0.0073687, 
    0.0073693, 0.0073694, 0.0073687, 0.0073682, 0.007368, 0.0073671, 
    0.007366, 0.0073646, 0.0073643, 0.0073651, 0.0073662, 0.0073671, 
    0.0073673, 0.0073675, 0.0073678, 0.0073674, 0.0073667, 0.0073647, 
    0.0073625, 0.0073599, 0.0073571, 0.0073543, 0.0073509, 0.0073471, 
    0.0073428, 0.0073384, 0.007334, 0.0073302, 0.0073272, 0.0073259, 
    0.0073257, 0.0073261, 0.0073262, 0.0073259, 0.0073246, 0.0073229, 
    0.0073211, 0.0073195, 0.0073181, 0.0073172, 0.0073166, 0.0073161, 
    0.0073144, 0.0073125, 0.0073103, 0.0073072, 0.0073035, 0.0072983, 
    0.0072928, 0.0072873, 0.0072818, 0.0072764, 0.0072715, 0.007267, 
    0.007264, 0.0072617, 0.0072603, 0.00726, 0.0072602, 0.0072612, 0.0072624, 
    0.0072636, 0.0072645, 0.0072652, 0.0072647, 0.007264, 0.0072627, 
    0.0072598, 0.0072562, 0.0072523, 0.0072485, 0.0072448, 0.0072415, 
    0.0072386, 0.0072361, 0.0072335, 0.0072306, 0.0072281, 0.007226, 
    0.0072238, 0.0072215, 0.0072187, 0.007216, 0.0072133, 0.0072105, 
    0.0072079, 0.0072058, 0.007203, 0.0071994, 0.0071959, 0.0071923, 
    0.0071883, 0.007184, 0.007179, 0.0071741, 0.007169, 0.0071634, 0.0071583, 
    0.0071539, 0.0071483, 0.0071422, 0.0071382, 0.0071341, 0.0071296, 
    0.0071247, 0.0071196, 0.0071145, 0.007109, 0.0071025, 0.0070954, 
    0.0070879, 0.0070805, 0.0070733, 0.0070664, 0.0070596, 0.0070527, 
    0.0070474, 0.0070425, 0.0070385, 0.0070348, 0.0070315, 0.0070284, 
    0.0070252, 0.0070216, 0.0070167, 0.0070103, 0.0070051, 0.0069999, 
    0.006994, 0.0069875, 0.0069804, 0.0069719, 0.0069628, 0.0069523, 
    0.0069416, 0.0069303, 0.0069189, 0.0069073, 0.0068951, 0.0068821, 
    0.0068674, 0.006853, 0.0068387, 0.0068246, 0.0068109, 0.006798, 
    0.0067868, 0.0067767, 0.0067659, 0.0067551, 0.0067442, 0.006733, 
    0.0067217, 0.0067103, 0.0066988, 0.0066869, 0.0066744, 0.0066613, 
    0.0066483, 0.0066354, 0.0066228, 0.0066111, 0.0066002, 0.0065915, 
    0.0065834, 0.0065755, 0.0065678, 0.0065604, 0.006555, 0.0065503, 
    0.0065468, 0.0065426, 0.0065372, 0.0065324, 0.0065279, 0.006525, 
    0.0065228, 0.0065218, 0.0065216, 0.0065218, 0.0065222, 0.0065224, 
    0.0065223, 0.0065223, 0.0065223, 0.0065228, 0.0065236, 0.0065249, 
    0.0065257, 0.0065262, 0.0065275, 0.0065288, 0.00653, 0.0065306, 
    0.0065308, 0.0065317, 0.0065324, 0.006531, 0.0065292, 0.0065268, 
    0.0065243, 0.0065216, 0.0065176, 0.0065134, 0.0065089, 0.006505, 
    0.0065012, 0.006497, 0.0064936, 0.0064911, 0.0064914, 0.0064927, 
    0.0064923, 0.0064915, 0.0064901, 0.006489, 0.006488, 0.0064869, 
    0.0064865, 0.0064875, 0.0064891, 0.006491, 0.0064907, 0.0064898, 
    0.0064872, 0.0064852, 0.0064835, 0.0064836, 0.006484, 0.0064852, 
    0.0064854, 0.0064848, 0.0064841, 0.0064838, 0.006485, 0.0064873, 
    0.0064908, 0.0064944, 0.0064982, 0.0065021, 0.0065062, 0.0065104, 
    0.0065146, 0.006519, 0.0065238, 0.0065286, 0.0065334, 0.0065377, 
    0.0065418, 0.0065458, 0.00655, 0.0065548, 0.0065591, 0.0065631, 
    0.0065679, 0.0065724, 0.0065763, 0.0065793, 0.0065817, 0.0065832, 
    0.0065845, 0.0065856, 0.0065873, 0.0065895, 0.0065896, 0.0065885, 
    0.0065841, 0.0065794, 0.0065744, 0.0065708, 0.0065673, 0.0065633, 
    0.0065589, 0.0065541, 0.0065501, 0.0065463, 0.0065425, 0.0065388, 
    0.0065353, 0.006532, 0.0065287, 0.0065245, 0.0065205, 0.0065165, 
    0.0065127, 0.0065091, 0.006504, 0.0064985, 0.0064921, 0.0064857, 
    0.0064791, 0.0064732, 0.0064675, 0.006462, 0.0064574, 0.0064533, 
    0.0064482, 0.0064433, 0.0064386, 0.0064348, 0.0064316, 0.006429, 
    0.0064266, 0.0064244, 0.0064229, 0.0064221, 0.0064214, 0.0064207, 
    0.0064201, 0.0064196, 0.0064193, 0.0064198, 0.0064204, 0.0064201, 
    0.0064195, 0.0064187, 0.0064178, 0.0064169, 0.0064161, 0.0064145, 
    0.0064117, 0.0064068, 0.0064009, 0.0063933, 0.0063857, 0.0063779, 
    0.0063699, 0.0063619, 0.0063537, 0.0063453, 0.0063363, 0.0063269, 
    0.0063172, 0.0063084, 0.0063003, 0.0062936, 0.0062883, 0.0062842, 
    0.0062803, 0.0062765, 0.0062725, 0.0062678, 0.0062626, 0.0062571, 
    0.0062516, 0.0062461, 0.0062405, 0.0062348, 0.0062287, 0.0062224, 
    0.0062147, 0.0062075, 0.0062006, 0.0061944, 0.0061885, 0.0061839, 
    0.0061803, 0.0061782, 0.0061781, 0.0061788, 0.0061813, 0.0061844, 
    0.0061884, 0.0061931, 0.0061981, 0.0062027, 0.0062065, 0.0062088, 
    0.0062101, 0.0062108, 0.0062111, 0.006211, 0.0062099, 0.006208, 
    0.0062053, 0.0062013, 0.0061969, 0.0061919, 0.0061865, 0.0061809, 
    0.0061775, 0.0061744, 0.0061713, 0.0061677, 0.0061637, 0.0061595, 
    0.0061552, 0.0061504, 0.0061457, 0.006141, 0.0061365, 0.0061319, 
    0.0061259, 0.006119, 0.0061106, 0.0061016, 0.0060922, 0.0060839, 
    0.0060759, 0.0060684, 0.0060615, 0.0060549, 0.0060492, 0.0060439, 
    0.0060395, 0.0060359, 0.0060329, 0.0060302, 0.0060276, 0.0060249, 
    0.0060213, 0.006017, 0.0060123, 0.0060075, 0.0060033, 0.0059991, 
    0.0059949, 0.0059913, 0.0059878, 0.0059843, 0.0059805, 0.0059766, 
    0.0059734, 0.0059704, 0.0059674, 0.0059647, 0.0059622, 0.0059586, 
    0.0059545, 0.0059501, 0.0059457, 0.0059412, 0.0059367, 0.0059322, 
    0.0059278, 0.0059225, 0.0059154, 0.0059073, 0.0058988, 0.0058886, 
    0.0058778, 0.0058657, 0.0058537, 0.0058416, 0.0058314, 0.0058219, 
    0.0058141, 0.005807, 0.0058004, 0.0057959, 0.0057917, 0.0057878, 
    0.0057839, 0.0057801, 0.0057767, 0.0057734, 0.0057695, 0.0057652, 
    0.0057605, 0.0057558, 0.0057511, 0.0057459, 0.0057404, 0.0057347, 
    0.0057289, 0.0057232, 0.005718, 0.0057129, 0.005708, 0.005703, 0.0056978, 
    0.0056919, 0.0056855, 0.0056779, 0.0056707, 0.0056636, 0.0056572, 
    0.005651, 0.0056456, 0.0056404, 0.0056354, 0.0056298, 0.0056241, 
    0.005618, 0.0056114, 0.0056042, 0.0055982, 0.0055922, 0.0055857, 
    0.0055792, 0.0055726, 0.0055658, 0.0055589, 0.0055522, 0.0055458, 
    0.0055397, 0.0055341, 0.0055287, 0.0055237, 0.0055188, 0.0055142, 
    0.0055094, 0.0055044, 0.0054991, 0.0054939, 0.0054889, 0.0054851, 
    0.0054819, 0.0054803, 0.0054793, 0.0054796, 0.0054801, 0.0054806, 
    0.0054825, 0.0054845, 0.0054866, 0.0054891, 0.0054919, 0.0054959, 
    0.0054999, 0.0055038, 0.0055067, 0.0055088, 0.0055098, 0.0055107, 
    0.005512, 0.0055133, 0.0055147, 0.0055159, 0.0055168, 0.0055162, 
    0.0055142, 0.0055107, 0.005507, 0.0055032, 0.0054994, 0.0054956, 
    0.0054918, 0.0054882, 0.0054847, 0.0054824, 0.0054804, 0.0054791, 
    0.005478, 0.0054769, 0.0054747, 0.0054724, 0.0054697, 0.005467, 
    0.0054643, 0.0054618, 0.0054591, 0.005456, 0.0054523, 0.0054484, 
    0.0054432, 0.0054375, 0.0054308, 0.0054247, 0.005419, 0.0054148, 
    0.0054105, 0.0054056, 0.0054003, 0.0053945, 0.0053882, 0.0053818, 
    0.0053755, 0.0053704, 0.0053667, 0.0053649, 0.0053636, 0.0053622, 
    0.0053605, 0.0053587, 0.0053567, 0.0053548, 0.0053527, 0.0053505, 
    0.0053482, 0.0053455, 0.0053426, 0.0053387, 0.0053345, 0.00533, 
    0.0053251, 0.00532, 0.0053142, 0.005308, 0.0053012, 0.0052939, 0.0052863, 
    0.0052796, 0.0052731, 0.0052668, 0.0052607, 0.0052548, 0.0052487, 
    0.0052425, 0.0052359, 0.0052292, 0.0052224, 0.0052152, 0.0052081, 
    0.0052017, 0.0051952, 0.0051887, 0.0051816, 0.0051744, 0.0051674, 
    0.0051608, 0.0051549, 0.0051501, 0.0051459, 0.0051427, 0.0051398, 
    0.0051373, 0.0051347, 0.0051323, 0.0051302, 0.0051282, 0.0051266, 
    0.0051249, 0.0051231, 0.0051213, 0.0051195, 0.005118, 0.0051161, 
    0.0051139, 0.0051121, 0.00511, 0.0051073, 0.0051047, 0.0051021, 
    0.0050995, 0.0050969, 0.0050946, 0.0050925, 0.0050906, 0.0050891, 
    0.0050877, 0.0050865, 0.0050852, 0.005084, 0.0050833, 0.0050828, 
    0.0050824, 0.005082, 0.0050815, 0.0050809, 0.0050801, 0.0050773, 
    0.0050741, 0.0050702, 0.0050665, 0.0050628, 0.0050582, 0.0050533, 
    0.0050478, 0.0050424, 0.0050373, 0.0050319, 0.0050267, 0.0050221, 
    0.0050183, 0.0050152, 0.0050129, 0.0050107, 0.0050083, 0.0050063, 
    0.0050045, 0.0050022, 0.0049996, 0.0049959, 0.0049919, 0.0049878, 
    0.0049831, 0.0049781, 0.0049722, 0.0049664, 0.0049607, 0.0049552, 
    0.0049498, 0.0049442, 0.0049389, 0.0049337, 0.0049284, 0.004923, 
    0.0049175, 0.0049123, 0.0049074, 0.0049029, 0.0048984, 0.0048939, 
    0.0048892, 0.0048839, 0.0048784, 0.0048728, 0.0048673, 0.0048624, 
    0.0048585, 0.0048544, 0.0048502, 0.004845, 0.0048398, 0.0048348, 
    0.0048295, 0.004824, 0.0048191, 0.0048144, 0.0048104, 0.0048071, 
    0.0048043, 0.0048016, 0.004799, 0.0047967, 0.0047948, 0.0047933, 
    0.0047921, 0.004791, 0.00479, 0.004789, 0.0047879, 0.0047859, 0.0047836, 
    0.0047809, 0.0047779, 0.0047745, 0.0047711, 0.0047677, 0.0047639, 
    0.0047602, 0.004757, 0.0047547, 0.0047529, 0.0047511, 0.0047493, 
    0.0047759, 0.004766, 0.0047561, 0.0047461, 0.0047361, 0.004726, 
    0.0047159, 0.0047058, 0.0046957, 0.0046856, 0.0046755, 0.0046654, 
    0.0046553, 0.0046454, 0.0046355, 0.0046256, 0.0046159, 0.0046062, 
    0.0045967, 0.0045873, 0.004578, 0.0045688, 0.0045597, 0.0045507, 
    0.0045418, 0.0045331, 0.0045244, 0.0045157, 0.0045072, 0.0044987, 
    0.0044902, 0.0044817, 0.0044732, 0.0044648, 0.0044563, 0.0044478, 
    0.0044392, 0.0044306, 0.004422, 0.0044133, 0.0044046, 0.0043959, 
    0.0043871, 0.0043783, 0.0043694, 0.0043606, 0.0043517, 0.0043428, 
    0.004334, 0.0043251, 0.0043163, 0.0043075, 0.0042987, 0.0042899, 
    0.0042812, 0.0042725, 0.0042639, 0.0042553, 0.0042467, 0.0042382, 
    0.0042297, 0.0042212, 0.0042127, 0.0042042, 0.0041957, 0.0041872, 
    0.0041787, 0.0041701, 0.0041615, 0.0041529, 0.0041442, 0.0041355, 
    0.0041267, 0.0041179, 0.004109, 0.0041001, 0.0040911, 0.0040821, 
    0.004073, 0.0040639, 0.0040548, 0.0040456, 0.0040364, 0.0040272, 
    0.004018, 0.0040088, 0.0039995, 0.0039903, 0.0039811, 0.0039719, 
    0.0039627, 0.0039535, 0.0039443, 0.0039352, 0.003926, 0.0039169, 
    0.0039078, 0.0038987, 0.0038896, 0.0038805, 0.0038714, 0.0038623, 
    0.0038532, 0.0038441, 0.0038351, 0.003826, 0.003817, 0.0038079, 
    0.0037988, 0.0037898, 0.0037807, 0.0037717, 0.0037626, 0.0037536, 
    0.0037445, 0.0037355, 0.0037264, 0.0037174, 0.0037083, 0.0036992, 
    0.0036902, 0.0036811, 0.003672, 0.003663, 0.0036539, 0.0036448, 
    0.0036357, 0.0036266, 0.0036175, 0.0036084, 0.0035993, 0.0035902, 
    0.0035811, 0.003572, 0.003563, 0.0035539, 0.0035448, 0.0035358, 
    0.0035267, 0.0035177, 0.0035087, 0.0034997, 0.0034908, 0.0034819, 
    0.003473, 0.0034642, 0.0034554, 0.0034467, 0.003438, 0.0034294, 
    0.0034208, 0.0034123, 0.0034039, 0.0033955, 0.0033871, 0.0033789, 
    0.0033706, 0.0033625, 0.0033543, 0.0033462, 0.0033382, 0.0033302, 
    0.0033222, 0.0033143, 0.0033064, 0.0032985, 0.0032907, 0.0032828, 
    0.003275, 0.0032672, 0.0032594, 0.0032517, 0.0032439, 0.0032361, 
    0.0032284, 0.0032206, 0.0032129, 0.0032051, 0.0031974, 0.0031896, 
    0.0031819, 0.0031741, 0.0031664, 0.0031586, 0.0031509, 0.0031431, 
    0.0031354, 0.0031276, 0.0031199, 0.0031121, 0.0031044, 0.0030966, 
    0.0030888, 0.0030811, 0.0030733, 0.0030655, 0.0030577, 0.0030499, 
    0.0030421, 0.0030343, 0.0030266, 0.0030188, 0.003011, 0.0030033, 
    0.0029956, 0.0029879, 0.0029802, 0.0029726, 0.0029651, 0.0029576, 
    0.0029502, 0.0029428, 0.0029355, 0.0029283, 0.0029211, 0.0029141, 
    0.0029071, 0.0029001, 0.0028933, 0.0028865, 0.0028797, 0.002873, 
    0.0028663, 0.0028597, 0.0028531, 0.0028465, 0.00284, 0.0028334, 
    0.0028269, 0.0028204, 0.0028138, 0.0028072, 0.0028006, 0.002794, 
    0.0027874, 0.0027808, 0.0027741, 0.0027674, 0.0027607, 0.002754, 
    0.0027472, 0.0027404, 0.0027337, 0.0027269, 0.00272, 0.0027132, 
    0.0027063, 0.0026994, 0.0026925, 0.0026856, 0.0026786, 0.0026716, 
    0.0026646, 0.0026575, 0.0026504, 0.0026432, 0.002636, 0.0026287, 
    0.0026214, 0.002614, 0.0026066, 0.002599, 0.0025915, 0.0025838, 
    0.0025761, 0.0025684, 0.0025606, 0.0025527, 0.0025448, 0.0025368, 
    0.0025288, 0.0025208, 0.0025128, 0.0025048, 0.0024967, 0.0024887, 
    0.0024807, 0.0024726, 0.0024647, 0.0024567, 0.0024488, 0.002441, 
    0.0024332, 0.0024254, 0.0024177, 0.00241, 0.0024024, 0.0023948, 
    0.0023873, 0.0023798, 0.0023723, 0.0023648, 0.0023574, 0.00235, 
    0.0023427, 0.0023353, 0.002328, 0.0023207, 0.0023134, 0.0023062, 
    0.0022989, 0.0022918, 0.0022846, 0.0022776, 0.0022706, 0.0022636, 
    0.0022567, 0.0022499, 0.0022431, 0.0022364, 0.0022298, 0.0022233, 
    0.0022168, 0.0022105, 0.0022042, 0.0021979, 0.0021918, 0.0021856, 
    0.0021796, 0.0021736, 0.0021677, 0.0021619, 0.002156, 0.0021503, 
    0.0021445, 0.0021389, 0.0021332, 0.0021276, 0.0021221, 0.0021165, 
    0.002111, 0.0021056, 0.0021001, 0.0020947, 0.0020892, 0.0020838, 
    0.0020784, 0.002073, 0.0020676, 0.0020622, 0.0020568, 0.0020513, 
    0.0020459, 0.0020404, 0.0020349, 0.0020294, 0.0020238, 0.0020182, 
    0.0020126, 0.0020069, 0.0020012, 0.0019955, 0.0019897, 0.0019839, 
    0.001978, 0.0019721, 0.0019662, 0.0019602, 0.0019542, 0.0019481, 
    0.0019419, 0.0019358, 0.0019296, 0.0019233, 0.001917, 0.0019107, 
    0.0019043, 0.0018979, 0.0018915, 0.001885, 0.0018785, 0.001872, 
    0.0018655, 0.0018589, 0.0018523, 0.0018457, 0.001839, 0.0018324, 
    0.0018257, 0.0018191, 0.0018124, 0.0018057, 0.001799, 0.0017924, 
    0.0017857, 0.001779, 0.0017723, 0.0017656, 0.001759, 0.0017523, 
    0.0017456, 0.0017389, 0.0017323, 0.0017256, 0.0017189, 0.0017123, 
    0.0017057, 0.001699, 0.0016924, 0.0016859, 0.0016793, 0.0016728, 
    0.0016663, 0.0016599, 0.0016535, 0.0016472, 0.001641, 0.0016348, 
    0.0016286, 0.0016226, 0.0016166, 0.0016106, 0.0016048, 0.001599, 
    0.0015932, 0.0015875, 0.0015819, 0.0015763, 0.0015707, 0.0015651, 
    0.0015596, 0.001554, 0.0015485, 0.0015429, 0.0015374, 0.0015318, 
    0.0015262, 0.0015206, 0.001515, 0.0015094, 0.0015037, 0.001498, 
    0.0014923, 0.0014865, 0.0014808, 0.001475, 0.0014692, 0.0014635, 
    0.0014577, 0.0014519, 0.0014462, 0.0014404, 0.0014347, 0.001429, 
    0.0014233, 0.0014176, 0.0014119, 0.0014063, 0.0014006, 0.001395, 
    0.0013894, 0.0013838, 0.0013782, 0.0013727, 0.0013671, 0.0013616, 
    0.001356, 0.0013505, 0.001345, 0.0013395, 0.001334, 0.0013286, 0.0013232, 
    0.0013179, 0.0013126, 0.0013073, 0.0013021, 0.001297, 0.0012919, 
    0.0012869, 0.0012819, 0.001277, 0.0012722, 0.0012675, 0.0012628, 
    0.0012581, 0.0012535, 0.001249, 0.0012444, 0.0012399, 0.0012355, 
    0.001231, 0.0012266, 0.0012222, 0.0012178, 0.0012133, 0.0012089, 
    0.0012044, 0.0011999, 0.0011954, 0.0011908, 0.0011862, 0.0011815, 
    0.0011768, 0.0011721, 0.0011672, 0.0011624, 0.0011574, 0.0011524, 
    0.0011474, 0.0011422, 0.0011371, 0.0011318, 0.0011265, 0.0011212, 
    0.0011158, 0.0011103, 0.0011049, 0.0010994, 0.0010939, 0.0010883, 
    0.0010828, 0.0010773, 0.0010719, 0.0010664, 0.0010611, 0.0010558, 
    0.0010505, 0.0010454, 0.0010403, 0.0010353, 0.0010304, 0.0010257, 
    0.001021, 0.0010164, 0.0010119, 0.0010076, 0.0010033, 0.00099918, 
    0.00099512, 0.00099115, 0.00098726, 0.00098344, 0.00097969, 0.000976, 
    0.00097236, 0.00096877, 0.00096521, 0.00096167, 0.00095816, 0.00095466, 
    0.00095116, 0.00094766, 0.00094416, 0.00094065, 0.00093712, 0.00093358, 
    0.00093002, 0.00092645, 0.00092286, 0.00091926, 0.00091565, 0.00091203, 
    0.00090841, 0.00090478, 0.00090115, 0.00089751, 0.00089388, 0.00089025, 
    0.00088661, 0.00088298, 0.00087933, 0.00087568, 0.00087202, 0.00086833, 
    0.00086462, 0.00086088, 0.00085711, 0.00085329, 0.00084943, 0.00084551, 
    0.00084155, 0.00083752, 0.00083344, 0.00082929, 0.00082509, 0.00082083, 
    0.00081653, 0.00081217, 0.00080777, 0.00080333, 0.00079887, 0.00079439, 
    0.00078989, 0.00078539, 0.00078089, 0.0007764, 0.00077194, 0.0007675, 
    0.00076309, 0.00075872, 0.0007544, 0.00075012, 0.00074589, 0.00074173, 
    0.00073761, 0.00073356, 0.00072958, 0.00072565, 0.0007218, 0.00071801, 
    0.0007143, 0.00071065, 0.00070708, 0.00070357, 0.00070015, 0.00069679, 
    0.00069351, 0.0006903, 0.00068716, 0.00068409, 0.00068108, 0.00067813, 
    0.00067523, 0.00067238, 0.00066957, 0.0006668, 0.00066406, 0.00066134, 
    0.00065863, 0.00065594, 0.00065325, 0.00065056, 0.00064788, 0.00064518, 
    0.00064248, 0.00063977, 0.00063704, 0.00063431, 0.00063157, 0.00062883, 
    0.00062607, 0.0006233, 0.00062052, 0.00061773, 0.00061494, 0.00061213, 
    0.00060931, 0.00060647, 0.00060363, 0.00060076, 0.00059788, 0.00059498, 
    0.00059206, 0.00058913, 0.00058618, 0.00058321, 0.00058023, 0.00057725, 
    0.00057425, 0.00057125, 0.00056825, 0.00056524, 0.00056224, 0.00055925, 
    0.00055625, 0.00055327, 0.00055028, 0.00054729, 0.00054431, 0.00054131, 
    0.0005383, 0.00053528, 0.00053224, 0.00052916, 0.00052606, 0.00052293, 
    0.00051976, 0.00051655, 0.0005133, 0.00051003, 0.00050672, 0.00050339, 
    0.00050004, 0.00049668, 0.00049332, 0.00048996, 0.00048662, 0.0004833, 
    0.00048001, 0.00047677, 0.00047357, 0.00047043, 0.00046735, 0.00046434, 
    0.0004614, 0.00045853, 0.00045574, 0.00045304, 0.00045042, 0.00044788, 
    0.00044544, 0.00044308, 0.0004408, 0.00043861, 0.00043651, 0.00043449, 
    0.00043256, 0.0004307, 0.00042891, 0.0004272, 0.00042555, 0.00042396, 
    0.00042242, 0.00042092, 0.00041946, 0.00041803, 0.00041661, 0.00041521, 
    0.00041381, 0.0004124, 0.00041098, 0.00040954, 0.00040807, 0.00040658, 
    0.00040505, 0.00040348, 0.00040186, 0.00040021, 0.00039851, 0.00039677, 
    0.00039499, 0.00039316, 0.00039129, 0.00038939, 0.00038745, 0.00038548, 
    0.00038347, 0.00038144, 0.00037938, 0.00037731, 0.0003752, 0.00037309, 
    0.00037096, 0.00036881, 0.00036666, 0.00036449, 0.00036232, 0.00036015, 
    0.00035798, 0.00035581, 0.00035364, 0.00035148, 0.00034932, 0.00034717, 
    0.00034503, 0.00034289, 0.00034077, 0.00033866, 0.00033655, 0.00033446, 
    0.00033238, 0.0003303, 0.00032824, 0.00032618, 0.00032413, 0.00032208, 
    0.00032004, 0.000318, 0.00031597, 0.00031394, 0.00031191, 0.00030988, 
    0.00030785, 0.00030582, 0.00030378, 0.00030174, 0.00029969, 0.00029763, 
    0.00029556, 0.00029348, 0.00029138, 0.00028928, 0.00028717, 0.00028504, 
    0.0002829, 0.00028076, 0.00027861, 0.00027646, 0.00027432, 0.00027218, 
    0.00027005, 0.00026794, 0.00026586, 0.0002638, 0.00026178, 0.00025979, 
    0.00025785, 0.00025596, 0.00025413, 0.00025234, 0.00025062, 0.00024895, 
    0.00024734, 0.00024579, 0.00024429, 0.00024285, 0.00024146, 0.00024012, 
    0.00023881, 0.00023755, 0.00023632, 0.00023511, 0.00023393, 0.00023277, 
    0.00023161, 0.00023047, 0.00022933, 0.00022818, 0.00022704, 0.00022588, 
    0.00022471, 0.00022353, 0.00022234, 0.00022113, 0.0002199, 0.00021866, 
    0.0002174, 0.00021612, 0.00021482, 0.00021351, 0.00021219, 0.00021085, 
    0.00020949, 0.00020813, 0.00020676, 0.00020538, 0.000204, 0.00020262, 
    0.00020124, 0.00019987, 0.0001985, 0.00019715, 0.00019581, 0.00019449, 
    0.00019318, 0.00019191, 0.00019066, 0.00018943, 0.00018824, 0.00018707, 
    0.00018594, 0.00018483, 0.00018376, 0.00018271, 0.00018168, 0.00018068, 
    0.0001797, 0.00017874, 0.00017779, 0.00017685, 0.00017592, 0.000175, 
    0.00017408, 0.00017317, 0.00017225, 0.00017134, 0.00017042, 0.0001695, 
    0.00016858, 0.00016767, 0.00016675, 0.00016584, 0.00016493, 0.00016403, 
    0.00016314, 0.00016226, 0.0001614, 0.00016054, 0.0001597, 0.00015888, 
    0.00015808, 0.00015729, 0.00015653, 0.00015578, 0.00015505, 0.00015433, 
    0.00015363, 0.00015295, 0.00015227, 0.00015161, 0.00015096, 0.00015031, 
    0.00014966, 0.00014902, 0.00014838, 0.00014773, 0.00014708, 0.00014642, 
    0.00014574, 0.00014506, 0.00014436, 0.00014364, 0.0001429, 0.00014215, 
    0.00014138, 0.00014058, 0.00013977, 0.00013894, 0.00013809, 0.00013722, 
    0.00013633, 0.00013544, 0.00013452, 0.0001336, 0.00013267, 0.00013172, 
    0.00013077, 0.00012982, 0.00012886, 0.0001279, 0.00012693, 0.00012596, 
    0.000125, 0.00012402, 0.00012306, 0.00012209, 0.00012113, 0.00012016, 
    0.00011921, 0.00011825, 0.00011731, 0.00011638, 0.00011546, 0.00011455, 
    0.00011366, 0.00011279, 0.00011194, 0.00011111, 0.00011031, 0.00010953, 
    0.00010879, 0.00010806, 0.00010737, 0.0001067, 0.00010605, 0.00010543, 
    0.00010483, 0.00010424, 0.00010366, 0.00010309, 0.00010253, 0.00010196, 
    0.00010139, 0.0001008, 0.00010021, 9.9604e-05, 9.8984e-05, 9.8344e-05, 
    9.7687e-05, 9.7018e-05, 9.6336e-05, 9.5646e-05, 9.4949e-05, 9.4252e-05, 
    9.3557e-05, 9.2871e-05, 9.2198e-05, 9.1542e-05, 9.0907e-05, 9.0301e-05, 
    8.9717e-05, 8.9172e-05, 8.8652e-05, 8.8171e-05, 8.7722e-05, 8.7307e-05, 
    8.6924e-05, 8.657e-05, 8.6249e-05, 8.5949e-05, 8.5672e-05, 8.5415e-05, 
    8.5172e-05, 8.4943e-05, 8.4717e-05, 8.4499e-05, 8.428e-05, 8.4056e-05, 
    8.3825e-05, 8.3583e-05, 8.3329e-05, 8.3054e-05, 8.2763e-05, 8.2447e-05, 
    8.2109e-05, 8.1744e-05, 8.1351e-05, 8.0928e-05, 8.0477e-05, 7.9994e-05, 
    7.9479e-05, 7.8936e-05, 7.8361e-05, 7.7758e-05, 7.7125e-05, 7.6466e-05, 
    7.5782e-05, 7.5075e-05, 7.4347e-05, 7.3605e-05, 7.2845e-05, 7.2074e-05, 
    7.13e-05, 7.0518e-05, 6.9739e-05, 6.896e-05, 6.8191e-05, 6.7433e-05, 
    6.669e-05, 6.5964e-05, 6.5259e-05, 6.4581e-05, 6.3929e-05, 6.3302e-05, 
    6.2713e-05, 6.2153e-05, 6.1629e-05, 6.1142e-05, 6.069e-05, 6.0278e-05, 
    5.99e-05, 5.9561e-05, 5.926e-05, 5.8993e-05, 5.8762e-05, 5.856e-05, 
    5.8389e-05, 5.8244e-05, 5.8127e-05, 5.803e-05, 5.7952e-05, 5.7886e-05, 
    5.7834e-05, 5.7788e-05, 5.7745e-05, 5.7707e-05, 5.7663e-05, 5.7616e-05, 
    5.7557e-05, 5.7493e-05, 5.7412e-05, 5.732e-05, 5.7211e-05, 5.7087e-05, 
    5.6946e-05, 5.679e-05, 5.6615e-05, 5.6426e-05, 5.6221e-05, 5.6002e-05, 
    5.577e-05, 5.5523e-05, 5.5263e-05, 5.4992e-05, 5.4711e-05, 5.4417e-05, 
    5.4114e-05, 5.3798e-05, 5.3475e-05, 5.3141e-05, 5.2795e-05, 5.2442e-05, 
    5.2076e-05, 5.1703e-05, 5.132e-05, 5.0927e-05, 5.0531e-05, 5.0123e-05, 
    4.9713e-05, 4.9297e-05, 4.8878e-05, 4.8457e-05, 4.8037e-05, 4.7619e-05, 
    4.7202e-05, 4.679e-05, 4.6384e-05, 4.5984e-05, 4.5589e-05, 4.5202e-05, 
    4.4823e-05, 4.4454e-05, 4.4089e-05, 4.3734e-05, 4.3386e-05, 4.3045e-05, 
    4.2709e-05, 4.2378e-05, 4.2057e-05, 4.1734e-05, 4.142e-05, 4.1108e-05, 
    4.08e-05, 4.0496e-05, 4.0198e-05, 3.9901e-05, 3.9611e-05, 3.9326e-05, 
    3.9047e-05, 3.8775e-05, 3.8512e-05, 3.8258e-05, 3.8011e-05, 3.7771e-05, 
    3.7546e-05, 3.7325e-05, 3.7112e-05, 3.6907e-05, 3.6708e-05, 3.6517e-05, 
    3.6327e-05, 3.6138e-05, 3.5954e-05, 3.5767e-05, 3.558e-05, 3.5391e-05, 
    3.5201e-05, 3.5003e-05, 3.4803e-05, 3.4598e-05, 3.4387e-05, 3.4175e-05, 
    3.3956e-05, 3.3733e-05, 3.3503e-05, 3.3271e-05, 3.3032e-05, 3.2792e-05, 
    3.2541e-05, 3.2287e-05, 3.2029e-05, 3.1766e-05, 3.1493e-05, 3.1217e-05, 
    3.0931e-05, 3.0643e-05, 3.0346e-05, 3.0046e-05, 2.9744e-05, 2.9437e-05, 
    2.9128e-05, 2.882e-05, 2.8514e-05, 2.8209e-05, 2.7909e-05, 2.7619e-05, 
    2.7335e-05, 2.7063e-05, 2.6798e-05, 2.6553e-05, 2.6315e-05, 2.6095e-05, 
    2.5892e-05, 2.57e-05, 2.5529e-05, 2.5366e-05, 2.5226e-05, 2.5094e-05, 
    2.498e-05, 2.4878e-05, 2.4783e-05, 2.4702e-05, 2.4629e-05, 2.4563e-05, 
    2.4503e-05, 2.445e-05, 2.4401e-05, 2.4352e-05, 2.4307e-05, 2.4266e-05, 
    2.422e-05, 2.4178e-05, 2.4135e-05, 2.4087e-05, 2.404e-05, 2.3985e-05, 
    2.3926e-05, 2.3867e-05, 2.3794e-05, 2.3713e-05, 2.363e-05, 2.3531e-05, 
    2.3424e-05, 2.3308e-05, 2.3179e-05, 2.3044e-05, 2.2901e-05, 2.2748e-05, 
    2.2597e-05, 2.2441e-05, 2.2288e-05, 2.214e-05, 2.2e-05, 2.1875e-05, 
    2.1769e-05, 2.1678e-05, 2.1616e-05, 2.1578e-05, 2.1576e-05, 2.1599e-05, 
    2.1656e-05, 2.1745e-05, 2.1869e-05, 2.2016e-05, 2.2196e-05, 2.2397e-05, 
    2.2611e-05, 2.2841e-05, 2.3074e-05, 2.3309e-05, 2.3536e-05, 2.3747e-05, 
    2.3934e-05, 2.4092e-05, 2.4215e-05, 2.4294e-05, 2.4331e-05, 2.431e-05, 
    2.4238e-05, 2.4109e-05, 2.3921e-05, 2.368e-05, 2.3378e-05, 2.3024e-05, 
    2.2621e-05, 2.2171e-05, 2.168e-05, 2.1161e-05, 2.0609e-05, 2.0042e-05, 
    1.9464e-05, 1.8879e-05, 1.83e-05, 1.7734e-05, 1.7183e-05, 1.6664e-05, 
    1.6171e-05, 1.5717e-05, 1.531e-05, 1.4943e-05, 1.4629e-05, 1.4364e-05, 
    1.4158e-05, 1.3999e-05, 1.3895e-05, 1.3846e-05, 1.3843e-05, 1.3891e-05, 
    1.3983e-05, 1.4116e-05, 1.429e-05, 1.4493e-05, 1.4724e-05, 1.4986e-05, 
    1.5264e-05, 1.5559e-05, 1.586e-05, 1.6173e-05, 1.6484e-05, 1.679e-05, 
    1.7087e-05, 1.7376e-05, 1.7642e-05, 1.7887e-05, 1.8107e-05, 1.8298e-05, 
    1.8451e-05, 1.8571e-05, 1.8649e-05, 1.8688e-05, 1.8682e-05, 1.8633e-05, 
    1.8541e-05, 1.8402e-05, 1.8223e-05, 1.8004e-05, 1.7747e-05, 1.7458e-05, 
    1.7135e-05, 1.6785e-05, 1.6419e-05, 1.603e-05, 1.5629e-05, 1.5218e-05, 
    1.4804e-05, 1.4383e-05, 1.3968e-05, 1.3557e-05, 1.3149e-05, 1.2754e-05, 
    1.2366e-05, 1.1991e-05, 1.1625e-05, 1.1269e-05, 1.0927e-05, 1.0596e-05, 
    1.0272e-05, 9.9654e-06, 9.6633e-06, 9.3721e-06, 9.0905e-06, 8.8216e-06, 
    8.5618e-06, 8.3137e-06, 8.0787e-06, 7.8568e-06, 7.6552e-06, 7.4652e-06, 
    7.2993e-06, 7.1575e-06, 7.0376e-06, 6.9454e-06, 6.8832e-06, 6.8563e-06, 
    6.8566e-06, 6.8922e-06, 6.9634e-06, 7.0669e-06, 7.203e-06, 7.3721e-06, 
    7.5704e-06, 7.7961e-06, 8.0403e-06, 8.3074e-06, 8.5888e-06, 8.8822e-06, 
    9.1807e-06, 9.4822e-06, 9.7829e-06, 1.0077e-05, 1.0363e-05, 1.0641e-05, 
    1.0898e-05, 1.114e-05, 1.1371e-05, 1.1579e-05, 1.1771e-05, 1.1947e-05, 
    1.2103e-05, 1.2244e-05, 1.2372e-05, 1.2489e-05, 1.2593e-05, 1.2689e-05, 
    1.2777e-05, 1.2859e-05, 1.294e-05, 1.3014e-05, 1.3092e-05, 1.3163e-05, 
    1.3236e-05, 1.3304e-05, 1.3374e-05, 1.3436e-05, 1.3497e-05, 1.3548e-05, 
    1.3594e-05, 1.3626e-05, 1.3647e-05, 1.3654e-05, 1.3644e-05, 1.3615e-05, 
    1.3572e-05, 1.3506e-05, 1.3419e-05, 1.3319e-05, 1.3197e-05, 1.3057e-05, 
    1.2905e-05, 1.2737e-05, 1.2565e-05, 1.2381e-05, 1.2196e-05, 1.2007e-05, 
    1.1824e-05, 1.1644e-05, 1.1468e-05, 1.1304e-05, 1.1149e-05, 1.1002e-05, 
    1.087e-05, 1.0744e-05, 1.0628e-05, 1.0516e-05, 1.041e-05, 1.0308e-05, 
    1.02e-05, 1.0091e-05, 9.974e-06, 9.8469e-06, 9.7105e-06, 9.5631e-06, 
    9.3933e-06, 9.216e-06, 9.0185e-06, 8.8077e-06, 8.5847e-06, 8.3473e-06, 
    8.1025e-06, 7.8502e-06, 7.5941e-06, 7.3353e-06, 7.0782e-06, 6.8269e-06, 
    6.5838e-06, 6.3511e-06, 6.128e-06, 5.9187e-06, 5.7272e-06, 5.5458e-06, 
    5.3817e-06, 5.2366e-06, 5.097e-06, 4.9778e-06, 4.8702e-06, 4.7685e-06, 
    4.6809e-06, 4.5996e-06, 4.529e-06, 4.4633e-06, 4.4084e-06, 4.3584e-06, 
    4.319e-06, 4.2896e-06, 4.2671e-06, 4.2625e-06, 4.2708e-06, 4.2936e-06, 
    4.3302e-06, 4.39e-06, 4.4642e-06, 4.5599e-06, 4.668e-06, 4.7949e-06, 
    4.9339e-06, 5.0876e-06, 5.2469e-06, 5.413e-06, 5.5809e-06, 5.7475e-06, 
    5.9056e-06, 6.059e-06, 6.1961e-06, 6.3213e-06, 6.4302e-06, 6.519e-06, 
    6.5893e-06, 6.6406e-06, 6.6732e-06, 6.6881e-06, 6.6855e-06, 6.6687e-06, 
    6.6363e-06, 6.5943e-06, 6.5444e-06, 6.4873e-06, 6.4251e-06, 6.3594e-06, 
    6.2931e-06, 6.2273e-06, 6.1615e-06, 6.0984e-06, 6.0387e-06, 5.9802e-06, 
    5.9276e-06, 5.8764e-06, 5.8275e-06, 5.7821e-06, 5.7392e-06, 5.6989e-06, 
    5.6587e-06, 5.6212e-06, 5.5812e-06, 5.5452e-06, 5.5071e-06, 5.4689e-06, 
    5.4304e-06, 5.3912e-06, 5.3526e-06, 5.3126e-06, 5.2709e-06, 5.232e-06, 
    5.1896e-06, 5.1487e-06, 5.1066e-06, 5.0645e-06, 5.0241e-06, 4.9816e-06, 
    4.9405e-06, 4.8955e-06, 4.8496e-06, 4.8055e-06, 4.7585e-06, 4.7052e-06, 
    4.6506e-06, 4.5918e-06, 4.5267e-06, 4.4553e-06, 4.3791e-06, 4.2923e-06, 
    4.1994e-06, 4.0992e-06, 3.987e-06, 3.8675e-06, 3.7415e-06, 3.6083e-06, 
    3.4651e-06, 3.32e-06, 3.1699e-06, 3.0198e-06, 2.8708e-06, 2.7273e-06, 
    2.5907e-06, 2.4643e-06, 2.3532e-06, 2.258e-06, 2.1861e-06, 2.1376e-06, 
    2.1167e-06, 2.1245e-06, 2.1661e-06, 2.2394e-06, 2.3472e-06, 2.4855e-06, 
    2.6608e-06, 2.8628e-06, 3.0953e-06, 3.3502e-06, 3.6252e-06, 3.9159e-06, 
    4.2166e-06, 4.52e-06, 4.8247e-06, 5.1204e-06, 5.4048e-06, 5.6715e-06, 
    5.9162e-06, 6.1358e-06, 6.3245e-06, 6.4807e-06, 6.6047e-06, 6.6943e-06, 
    6.748e-06, 6.7684e-06, 6.756e-06, 6.7137e-06, 6.6421e-06, 6.5457e-06, 
    6.4269e-06, 6.2895e-06, 6.1369e-06, 5.9714e-06, 5.7971e-06, 5.6162e-06, 
    5.4322e-06, 5.247e-06, 5.0619e-06, 4.8802e-06, 4.701e-06, 4.527e-06, 
    4.3569e-06, 4.1916e-06, 4.0329e-06, 3.8764e-06, 3.7263e-06, 3.5792e-06, 
    3.4362e-06, 3.2962e-06, 3.1569e-06, 3.0218e-06, 2.8861e-06, 2.7542e-06, 
    2.6213e-06, 2.4898e-06, 2.3602e-06, 2.2309e-06, 2.1045e-06, 1.981e-06, 
    1.8572e-06, 1.7386e-06, 1.6236e-06, 1.5136e-06, 1.4095e-06, 1.312e-06, 
    1.2223e-06, 1.1404e-06, 1.0704e-06, 1.0096e-06, 9.6156e-07, 9.2663e-07, 
    9.0425e-07, 8.974e-07, 9.0491e-07, 9.2707e-07, 9.6319e-07, 1.0155e-06, 
    1.081e-06, 1.1618e-06, 1.2556e-06, 1.3615e-06, 1.4797e-06, 1.608e-06, 
    1.7458e-06, 1.8942e-06, 2.0486e-06, 2.2119e-06, 2.3789e-06, 2.5515e-06 ;

 bangle_opt =
  0.016718, 0.016852, 0.017001, 0.017179, 0.01739, 0.017619, 0.017865, 
    0.018113, 0.018368, 0.018649, 0.018947, 0.019248, 0.019549, 0.019851, 
    0.020152, 0.020453, 0.020723, 0.020983, 0.021224, 0.02145, 0.021662, 
    0.021837, 0.021995, 0.0221, 0.022208, 0.022319, 0.022431, 0.022541, 
    0.022629, 0.022716, 0.022803, 0.022899, 0.022999, 0.023103, 0.023203, 
    0.023296, 0.023372, 0.023442, 0.023487, 0.023527, 0.023554, 0.023578, 
    0.0236, 0.023595, 0.023582, 0.023553, 0.023522, 0.023488, 0.023466, 
    0.023443, 0.02342, 0.023396, 0.023372, 0.023346, 0.023321, 0.023301, 
    0.023285, 0.023273, 0.023284, 0.0233, 0.023316, 0.02333, 0.023342, 
    0.023331, 0.023312, 0.023286, 0.023263, 0.023245, 0.023228, 0.023209, 
    0.02318, 0.023147, 0.023109, 0.02308, 0.023055, 0.023048, 0.023045, 
    0.023048, 0.02305, 0.02305, 0.023051, 0.02306, 0.023089, 0.023127, 
    0.023171, 0.023203, 0.023232, 0.023259, 0.023284, 0.023309, 0.023337, 
    0.023366, 0.023397, 0.023423, 0.023444, 0.023459, 0.023473, 0.023483, 
    0.023494, 0.023503, 0.023507, 0.02351, 0.023515, 0.023519, 0.023525, 
    0.023529, 0.023533, 0.023531, 0.023526, 0.023517, 0.023513, 0.023511, 
    0.02351, 0.023505, 0.023493, 0.023478, 0.023462, 0.023443, 0.023423, 
    0.023401, 0.02338, 0.023361, 0.023351, 0.023342, 0.023334, 0.023327, 
    0.023321, 0.023327, 0.023334, 0.023341, 0.023349, 0.023356, 0.02337, 
    0.023386, 0.023405, 0.023423, 0.023441, 0.02346, 0.023478, 0.023492, 
    0.023507, 0.023522, 0.02354, 0.023559, 0.023574, 0.023591, 0.023611, 
    0.023635, 0.02366, 0.023686, 0.02371, 0.02373, 0.023763, 0.023803, 
    0.023851, 0.023897, 0.023934, 0.023982, 0.024036, 0.024096, 0.024154, 
    0.024207, 0.024256, 0.024302, 0.024348, 0.024393, 0.024436, 0.024479, 
    0.024522, 0.024568, 0.024614, 0.024652, 0.024688, 0.024724, 0.024762, 
    0.024802, 0.024846, 0.024894, 0.024949, 0.025003, 0.025057, 0.025111, 
    0.025169, 0.025233, 0.025298, 0.025364, 0.025408, 0.025446, 0.025476, 
    0.025487, 0.025489, 0.025428, 0.02535, 0.025231, 0.025113, 0.024996, 
    0.024862, 0.024724, 0.024574, 0.024431, 0.024294, 0.024187, 0.024083, 
    0.023971, 0.023857, 0.023742, 0.023623, 0.023499, 0.023352, 0.023204, 
    0.023055, 0.022906, 0.022753, 0.022574, 0.022377, 0.022156, 0.021965, 
    0.021785, 0.021608, 0.021428, 0.021245, 0.021053, 0.020858, 0.020655, 
    0.020456, 0.020267, 0.020092, 0.019925, 0.019811, 0.019708, 0.019628, 
    0.019582, 0.019559, 0.019539, 0.019518, 0.019494, 0.019472, 0.019451, 
    0.019406, 0.019349, 0.019258, 0.01916, 0.019055, 0.01897, 0.018886, 
    0.018788, 0.018696, 0.018611, 0.018527, 0.018442, 0.01834, 0.018264, 
    0.018223, 0.018205, 0.018191, 0.018136, 0.01807, 0.017985, 0.017913, 
    0.017847, 0.017749, 0.017665, 0.017611, 0.017562, 0.017516, 0.017454, 
    0.017394, 0.01734, 0.017289, 0.017242, 0.017195, 0.01715, 0.017109, 
    0.01707, 0.017032, 0.016995, 0.016962, 0.016949, 0.016947, 0.016957, 
    0.016973, 0.016987, 0.016989, 0.017005, 0.017039, 0.017079, 0.017121, 
    0.017168, 0.017217, 0.017269, 0.017302, 0.017328, 0.017347, 0.017371, 
    0.017402, 0.017449, 0.017503, 0.017545, 0.0176, 0.017679, 0.017726, 
    0.017755, 0.017787, 0.017814, 0.017827, 0.017834, 0.017837, 0.017837, 
    0.017836, 0.017827, 0.017817, 0.017807, 0.017794, 0.017781, 0.017769, 
    0.017757, 0.017744, 0.017734, 0.017727, 0.017729, 0.017737, 0.017749, 
    0.017752, 0.017752, 0.017742, 0.017728, 0.017711, 0.017677, 0.017637, 
    0.017594, 0.017551, 0.01751, 0.017471, 0.017432, 0.017394, 0.017357, 
    0.017321, 0.01729, 0.017263, 0.017244, 0.017233, 0.017237, 0.017259, 
    0.017291, 0.017329, 0.017369, 0.01741, 0.017451, 0.017492, 0.017539, 
    0.017585, 0.017629, 0.017668, 0.017704, 0.017737, 0.017767, 0.017789, 
    0.017805, 0.017815, 0.017822, 0.017828, 0.017842, 0.017856, 0.017871, 
    0.017902, 0.01794, 0.017996, 0.01805, 0.018102, 0.01815, 0.018195, 
    0.018238, 0.018281, 0.018322, 0.01836, 0.018397, 0.018428, 0.018458, 
    0.018482, 0.018496, 0.018502, 0.018502, 0.018501, 0.0185, 0.018499, 
    0.018497, 0.018495, 0.018491, 0.018485, 0.018482, 0.018481, 0.018481, 
    0.018482, 0.018482, 0.018481, 0.018477, 0.018463, 0.018448, 0.018429, 
    0.018411, 0.018391, 0.018371, 0.018351, 0.018332, 0.018313, 0.018295, 
    0.018276, 0.018256, 0.018242, 0.018231, 0.018222, 0.018211, 0.018198, 
    0.018197, 0.018196, 0.018198, 0.018193, 0.018184, 0.018175, 0.018167, 
    0.018161, 0.018154, 0.018146, 0.018136, 0.018125, 0.018118, 0.018111, 
    0.018105, 0.018097, 0.018089, 0.018086, 0.018085, 0.018086, 0.018087, 
    0.018089, 0.018095, 0.018104, 0.018116, 0.018127, 0.018136, 0.018139, 
    0.018138, 0.018131, 0.018124, 0.018117, 0.018114, 0.018111, 0.018105, 
    0.018097, 0.018086, 0.018081, 0.018073, 0.018059, 0.018047, 0.018035, 
    0.018037, 0.018039, 0.018038, 0.018032, 0.018024, 0.018027, 0.018032, 
    0.018041, 0.018044, 0.018042, 0.018034, 0.018024, 0.018017, 0.018007, 
    0.017994, 0.017986, 0.017978, 0.017972, 0.017963, 0.017951, 0.017944, 
    0.017937, 0.017938, 0.017943, 0.017954, 0.017972, 0.017994, 0.018011, 
    0.018029, 0.018047, 0.018067, 0.018088, 0.018106, 0.018122, 0.018132, 
    0.018139, 0.018146, 0.018151, 0.018155, 0.018154, 0.018154, 0.018156, 
    0.018156, 0.018154, 0.018144, 0.018135, 0.018127, 0.018129, 0.018133, 
    0.018138, 0.018143, 0.018147, 0.018152, 0.018157, 0.018159, 0.018164, 
    0.018171, 0.018178, 0.018184, 0.018183, 0.01818, 0.018177, 0.018171, 
    0.018163, 0.018156, 0.018149, 0.018143, 0.018134, 0.018124, 0.018111, 
    0.018099, 0.018091, 0.018087, 0.018085, 0.018082, 0.018078, 0.018073, 
    0.018068, 0.018064, 0.01806, 0.018056, 0.018053, 0.018049, 0.018044, 
    0.018036, 0.018028, 0.018019, 0.018011, 0.018003, 0.017995, 0.017986, 
    0.017979, 0.017971, 0.017963, 0.017955, 0.017948, 0.017941, 0.017934, 
    0.017927, 0.017921, 0.017914, 0.017908, 0.017901, 0.017895, 0.017891, 
    0.017888, 0.017885, 0.017881, 0.017877, 0.017875, 0.017874, 0.017876, 
    0.017879, 0.017883, 0.017888, 0.017893, 0.017897, 0.017901, 0.017905, 
    0.017908, 0.017912, 0.017918, 0.017924, 0.01793, 0.017931, 0.017926, 
    0.01792, 0.017913, 0.017911, 0.017906, 0.017898, 0.017889, 0.01788, 
    0.01787, 0.01786, 0.01785, 0.017839, 0.017827, 0.017816, 0.017805, 
    0.017795, 0.017785, 0.017775, 0.017761, 0.017749, 0.017737, 0.017725, 
    0.017712, 0.017696, 0.017679, 0.01766, 0.017639, 0.017615, 0.017592, 
    0.017569, 0.017545, 0.017522, 0.0175, 0.01748, 0.017461, 0.017443, 
    0.017427, 0.017414, 0.017408, 0.017403, 0.017396, 0.017389, 0.017379, 
    0.017375, 0.017373, 0.017372, 0.017371, 0.01737, 0.017369, 0.017369, 
    0.017368, 0.017367, 0.017365, 0.017363, 0.01736, 0.017354, 0.017347, 
    0.017336, 0.017323, 0.01731, 0.017297, 0.017284, 0.017272, 0.01726, 
    0.01725, 0.017243, 0.017236, 0.017231, 0.017227, 0.017223, 0.017221, 
    0.017218, 0.017214, 0.01721, 0.017208, 0.017206, 0.017205, 0.017206, 
    0.017208, 0.017211, 0.017212, 0.017213, 0.017211, 0.017209, 0.017208, 
    0.017208, 0.017208, 0.017208, 0.017209, 0.017209, 0.017205, 0.017198, 
    0.01719, 0.017186, 0.017188, 0.017191, 0.017195, 0.017204, 0.017215, 
    0.017232, 0.017251, 0.01727, 0.017291, 0.017312, 0.017332, 0.017353, 
    0.017373, 0.017394, 0.017416, 0.017436, 0.017454, 0.01747, 0.017482, 
    0.017492, 0.017497, 0.017501, 0.017502, 0.017504, 0.017507, 0.017507, 
    0.017506, 0.017501, 0.017492, 0.017481, 0.017467, 0.017453, 0.017438, 
    0.017424, 0.017412, 0.017407, 0.017402, 0.017396, 0.017387, 0.017377, 
    0.01737, 0.017364, 0.017357, 0.017347, 0.017335, 0.017323, 0.017312, 
    0.017304, 0.017294, 0.017284, 0.017272, 0.017259, 0.017246, 0.017233, 
    0.017221, 0.017209, 0.017199, 0.017191, 0.017185, 0.01718, 0.017177, 
    0.017174, 0.017168, 0.017163, 0.01716, 0.017158, 0.017156, 0.017157, 
    0.017161, 0.017169, 0.017177, 0.017187, 0.017196, 0.017205, 0.017213, 
    0.017222, 0.017231, 0.017244, 0.017257, 0.01727, 0.017282, 0.017293, 
    0.017304, 0.017317, 0.017332, 0.017347, 0.017362, 0.017381, 0.017402, 
    0.017433, 0.017466, 0.017501, 0.017538, 0.017577, 0.017625, 0.017674, 
    0.017723, 0.017771, 0.017819, 0.017857, 0.017893, 0.017924, 0.017954, 
    0.017985, 0.018018, 0.018049, 0.018078, 0.018103, 0.018124, 0.018144, 
    0.018164, 0.018185, 0.018206, 0.018227, 0.018244, 0.01826, 0.018273, 
    0.018286, 0.018297, 0.018306, 0.018314, 0.01832, 0.018323, 0.018325, 
    0.018326, 0.018324, 0.018315, 0.018303, 0.018289, 0.018271, 0.01825, 
    0.018222, 0.01819, 0.018153, 0.018109, 0.018062, 0.018011, 0.017963, 
    0.017918, 0.017872, 0.017824, 0.017767, 0.01771, 0.017652, 0.017594, 
    0.017535, 0.017477, 0.017417, 0.017356, 0.017289, 0.017219, 0.017147, 
    0.017074, 0.016998, 0.016922, 0.016844, 0.016764, 0.016684, 0.016605, 
    0.016525, 0.016442, 0.016357, 0.016273, 0.016191, 0.016111, 0.016032, 
    0.015949, 0.015865, 0.015785, 0.015707, 0.015631, 0.015556, 0.015482, 
    0.015416, 0.015353, 0.015292, 0.015234, 0.015177, 0.015134, 0.015093, 
    0.01506, 0.015026, 0.014992, 0.01496, 0.014929, 0.014899, 0.01487, 
    0.014842, 0.014821, 0.014802, 0.014786, 0.014772, 0.01476, 0.014749, 
    0.01474, 0.014734, 0.014729, 0.014724, 0.014719, 0.014715, 0.014713, 
    0.01471, 0.014708, 0.014704, 0.0147, 0.014695, 0.014689, 0.014681, 
    0.014671, 0.014661, 0.014652, 0.014643, 0.014634, 0.014621, 0.014608, 
    0.014597, 0.014585, 0.014569, 0.014551, 0.014532, 0.014518, 0.014503, 
    0.014488, 0.014472, 0.014456, 0.014443, 0.014431, 0.01442, 0.014409, 
    0.014398, 0.014385, 0.014372, 0.014357, 0.014343, 0.014328, 0.014315, 
    0.014303, 0.01429, 0.014275, 0.014258, 0.014239, 0.01422, 0.014203, 
    0.014186, 0.014169, 0.014153, 0.014138, 0.014122, 0.014105, 0.014086, 
    0.01407, 0.014056, 0.014046, 0.014035, 0.014024, 0.014016, 0.014009, 
    0.014001, 0.013993, 0.013986, 0.013981, 0.013977, 0.013974, 0.01397, 
    0.013965, 0.013959, 0.013953, 0.013946, 0.01394, 0.013935, 0.01393, 
    0.013926, 0.013922, 0.013917, 0.013908, 0.013902, 0.013897, 0.013894, 
    0.013891, 0.013889, 0.013888, 0.013885, 0.013885, 0.013887, 0.013887, 
    0.013889, 0.013891, 0.013895, 0.013899, 0.013892, 0.013885, 0.013879, 
    0.013876, 0.013873, 0.013866, 0.013858, 0.013852, 0.013847, 0.013842, 
    0.013837, 0.013834, 0.013834, 0.013836, 0.013838, 0.01384, 0.013842, 
    0.013843, 0.013845, 0.013849, 0.013852, 0.013855, 0.013858, 0.013861, 
    0.013864, 0.013865, 0.013866, 0.013866, 0.013867, 0.013869, 0.013871, 
    0.013873, 0.013874, 0.013874, 0.013875, 0.013875, 0.013875, 0.013876, 
    0.013879, 0.013886, 0.013891, 0.013895, 0.013896, 0.013899, 0.013905, 
    0.013909, 0.01391, 0.013913, 0.013915, 0.013917, 0.013917, 0.013914, 
    0.01391, 0.013906, 0.013902, 0.013899, 0.013896, 0.013892, 0.013886, 
    0.013876, 0.013865, 0.013853, 0.013842, 0.013831, 0.01382, 0.01381, 
    0.0138, 0.013789, 0.013778, 0.013765, 0.013754, 0.013744, 0.013736, 
    0.013729, 0.013719, 0.013711, 0.013704, 0.013695, 0.013686, 0.013679, 
    0.013672, 0.013664, 0.013655, 0.013647, 0.013637, 0.013626, 0.013616, 
    0.013606, 0.013594, 0.013582, 0.01357, 0.013559, 0.013547, 0.013535, 
    0.013524, 0.013513, 0.013502, 0.013495, 0.013491, 0.013487, 0.013482, 
    0.013483, 0.013482, 0.013479, 0.01348, 0.013481, 0.013483, 0.013484, 
    0.013481, 0.013477, 0.013471, 0.013466, 0.013461, 0.013459, 0.013455, 
    0.01345, 0.013447, 0.013443, 0.013438, 0.013432, 0.013427, 0.013424, 
    0.013423, 0.013428, 0.013429, 0.013429, 0.013428, 0.013427, 0.013428, 
    0.013429, 0.013429, 0.013429, 0.013429, 0.01343, 0.013431, 0.013432, 
    0.01343, 0.013428, 0.01343, 0.01343, 0.013429, 0.013431, 0.013434, 
    0.013427, 0.013422, 0.013418, 0.013418, 0.013418, 0.013417, 0.013415, 
    0.013411, 0.013405, 0.013397, 0.01339, 0.013383, 0.013374, 0.013367, 
    0.01336, 0.013355, 0.013348, 0.013339, 0.013329, 0.013317, 0.013308, 
    0.013299, 0.013289, 0.013277, 0.013266, 0.013256, 0.013246, 0.013237, 
    0.013227, 0.013217, 0.013205, 0.013193, 0.013183, 0.013171, 0.013157, 
    0.013144, 0.01313, 0.013114, 0.013101, 0.013092, 0.013081, 0.013068, 
    0.013057, 0.013046, 0.013036, 0.013028, 0.013022, 0.013017, 0.013013, 
    0.01301, 0.013007, 0.013005, 0.013, 0.012995, 0.01299, 0.012985, 0.01298, 
    0.012975, 0.012971, 0.012966, 0.012964, 0.012962, 0.01296, 0.012957, 
    0.012956, 0.012954, 0.012951, 0.012949, 0.012947, 0.012947, 0.012949, 
    0.012951, 0.012952, 0.012952, 0.012953, 0.012955, 0.012956, 0.012957, 
    0.012958, 0.012961, 0.012963, 0.012967, 0.012971, 0.012977, 0.012977, 
    0.012977, 0.012978, 0.012977, 0.012973, 0.012969, 0.012964, 0.01296, 
    0.012957, 0.012955, 0.012952, 0.012949, 0.012945, 0.012941, 0.012936, 
    0.012931, 0.012927, 0.012924, 0.012921, 0.012918, 0.012916, 0.012913, 
    0.012908, 0.012904, 0.0129, 0.012896, 0.012893, 0.012888, 0.012884, 
    0.012882, 0.01288, 0.012878, 0.012875, 0.012872, 0.012866, 0.012857, 
    0.012846, 0.012837, 0.012829, 0.012823, 0.012814, 0.012805, 0.012794, 
    0.012785, 0.012778, 0.01277, 0.012763, 0.012753, 0.012744, 0.012739, 
    0.012734, 0.01273, 0.012726, 0.012722, 0.012718, 0.012712, 0.012705, 
    0.012697, 0.012689, 0.012683, 0.012679, 0.012676, 0.01267, 0.012663, 
    0.012657, 0.012651, 0.012646, 0.012639, 0.012631, 0.012623, 0.012615, 
    0.012607, 0.012602, 0.012599, 0.012597, 0.012596, 0.012596, 0.012595, 
    0.012594, 0.012597, 0.012601, 0.012607, 0.012612, 0.012617, 0.012621, 
    0.012625, 0.012628, 0.01263, 0.012631, 0.012633, 0.012634, 0.012635, 
    0.012636, 0.012638, 0.01264, 0.012643, 0.012645, 0.012648, 0.012651, 
    0.012652, 0.012652, 0.01265, 0.012648, 0.012646, 0.012644, 0.012642, 
    0.012639, 0.012636, 0.012633, 0.012629, 0.012625, 0.01262, 0.012616, 
    0.012611, 0.012607, 0.012602, 0.012596, 0.01259, 0.012584, 0.012579, 
    0.012573, 0.012569, 0.012564, 0.01256, 0.012555, 0.012551, 0.012546, 
    0.01254, 0.012534, 0.012527, 0.012519, 0.012511, 0.012503, 0.012496, 
    0.012487, 0.012477, 0.012467, 0.012457, 0.012452, 0.012447, 0.012443, 
    0.01244, 0.012437, 0.012435, 0.012432, 0.012428, 0.012424, 0.012419, 
    0.012415, 0.012411, 0.012406, 0.012399, 0.012391, 0.012381, 0.012373, 
    0.012366, 0.01236, 0.012355, 0.012348, 0.012341, 0.012335, 0.01233, 
    0.012325, 0.01232, 0.012314, 0.012309, 0.012306, 0.012304, 0.0123, 
    0.012295, 0.01229, 0.012286, 0.012283, 0.012279, 0.012275, 0.012273, 
    0.012271, 0.012269, 0.012267, 0.012264, 0.012256, 0.012249, 0.012245, 
    0.012241, 0.012237, 0.012232, 0.012226, 0.012218, 0.012211, 0.012206, 
    0.012204, 0.012203, 0.012203, 0.012201, 0.012198, 0.012191, 0.012185, 
    0.012181, 0.012176, 0.01217, 0.012165, 0.012159, 0.012153, 0.012147, 
    0.012139, 0.012131, 0.012124, 0.012119, 0.012114, 0.012108, 0.012101, 
    0.012093, 0.012088, 0.012081, 0.012071, 0.012058, 0.012043, 0.012031, 
    0.01202, 0.01201, 0.012, 0.011988, 0.011977, 0.011967, 0.011959, 
    0.011951, 0.011942, 0.011934, 0.011925, 0.011917, 0.011908, 0.011898, 
    0.011888, 0.011878, 0.011868, 0.011859, 0.01185, 0.01184, 0.01183, 
    0.011821, 0.011813, 0.011806, 0.011799, 0.011792, 0.011784, 0.011778, 
    0.011773, 0.011768, 0.011764, 0.01176, 0.011755, 0.01175, 0.011747, 
    0.011746, 0.011745, 0.011745, 0.011744, 0.011743, 0.01174, 0.011738, 
    0.011736, 0.011735, 0.011735, 0.011735, 0.011734, 0.011733, 0.01173, 
    0.011726, 0.011723, 0.011721, 0.011721, 0.011723, 0.011723, 0.011721, 
    0.01172, 0.011719, 0.011717, 0.011715, 0.011714, 0.011711, 0.011708, 
    0.011707, 0.011706, 0.011705, 0.011702, 0.011698, 0.011694, 0.011691, 
    0.011687, 0.011681, 0.011675, 0.01167, 0.011666, 0.011663, 0.011658, 
    0.011652, 0.011647, 0.011642, 0.011639, 0.011636, 0.011633, 0.011629, 
    0.011625, 0.011622, 0.011619, 0.011616, 0.01161, 0.011605, 0.011602, 
    0.011598, 0.011592, 0.011589, 0.011586, 0.011581, 0.011577, 0.011574, 
    0.011572, 0.01157, 0.011569, 0.011567, 0.011565, 0.011564, 0.011563, 
    0.01156, 0.011558, 0.011556, 0.011554, 0.011554, 0.011553, 0.011552, 
    0.011551, 0.011549, 0.011546, 0.011544, 0.011542, 0.01154, 0.011538, 
    0.011535, 0.011529, 0.011524, 0.011519, 0.011514, 0.01151, 0.011506, 
    0.011501, 0.011497, 0.011492, 0.011486, 0.011478, 0.011471, 0.011465, 
    0.01146, 0.011457, 0.011451, 0.011445, 0.011438, 0.011431, 0.011424, 
    0.011415, 0.011406, 0.011397, 0.01139, 0.011385, 0.01138, 0.011376, 
    0.011371, 0.011365, 0.01136, 0.011356, 0.011351, 0.011348, 0.011345, 
    0.011344, 0.011341, 0.011338, 0.011335, 0.011332, 0.011328, 0.011324, 
    0.011319, 0.011314, 0.011309, 0.011303, 0.011297, 0.011292, 0.011289, 
    0.011286, 0.011285, 0.011283, 0.011281, 0.011276, 0.011272, 0.011269, 
    0.011267, 0.011266, 0.011267, 0.011268, 0.011268, 0.011267, 0.011265, 
    0.011262, 0.011258, 0.011254, 0.011251, 0.011247, 0.011244, 0.01124, 
    0.011237, 0.011233, 0.011228, 0.011224, 0.011219, 0.011215, 0.011211, 
    0.011208, 0.011205, 0.011203, 0.011204, 0.011204, 0.011204, 0.011203, 
    0.011202, 0.011199, 0.011195, 0.011194, 0.011192, 0.011192, 0.011191, 
    0.01119, 0.011189, 0.011187, 0.011184, 0.011181, 0.011178, 0.011174, 
    0.011171, 0.011169, 0.011167, 0.011165, 0.011161, 0.011158, 0.011154, 
    0.011151, 0.011148, 0.011142, 0.011137, 0.011135, 0.011135, 0.011135, 
    0.011135, 0.011134, 0.011133, 0.011132, 0.011131, 0.011129, 0.011127, 
    0.011125, 0.011123, 0.011122, 0.011124, 0.011125, 0.011127, 0.011128, 
    0.011126, 0.011124, 0.011121, 0.01112, 0.011121, 0.011122, 0.011122, 
    0.011121, 0.011119, 0.011117, 0.011113, 0.01111, 0.011108, 0.011105, 
    0.011103, 0.011101, 0.011098, 0.011095, 0.01109, 0.011086, 0.011082, 
    0.011075, 0.011067, 0.011061, 0.011055, 0.011051, 0.011047, 0.011043, 
    0.01104, 0.011037, 0.011032, 0.011027, 0.01102, 0.011016, 0.011012, 
    0.011008, 0.011002, 0.010995, 0.010989, 0.010982, 0.010976, 0.010968, 
    0.01096, 0.010951, 0.010942, 0.010934, 0.010926, 0.010918, 0.010911, 
    0.010903, 0.010895, 0.010888, 0.010881, 0.010875, 0.01087, 0.010864, 
    0.010858, 0.010854, 0.010851, 0.010849, 0.010845, 0.010842, 0.010837, 
    0.010831, 0.010824, 0.010819, 0.010812, 0.010804, 0.010798, 0.010794, 
    0.010788, 0.010783, 0.010775, 0.010768, 0.010761, 0.010756, 0.010752, 
    0.010748, 0.010745, 0.010741, 0.01074, 0.010739, 0.010737, 0.010736, 
    0.010735, 0.010734, 0.010734, 0.010735, 0.010737, 0.010738, 0.010737, 
    0.010735, 0.010731, 0.010727, 0.010725, 0.010722, 0.010721, 0.010719, 
    0.010716, 0.010709, 0.010702, 0.010696, 0.010692, 0.01069, 0.010692, 
    0.010695, 0.010697, 0.010696, 0.010694, 0.010693, 0.010691, 0.010689, 
    0.01069, 0.010691, 0.010691, 0.010691, 0.01069, 0.010687, 0.010684, 
    0.01068, 0.010676, 0.010673, 0.01067, 0.010668, 0.010663, 0.010658, 
    0.010653, 0.010647, 0.010642, 0.010641, 0.01064, 0.010641, 0.010641, 
    0.010641, 0.010637, 0.010633, 0.010631, 0.010631, 0.010632, 0.010634, 
    0.010635, 0.010633, 0.010628, 0.010618, 0.010612, 0.010607, 0.010603, 
    0.0106, 0.010599, 0.010596, 0.010591, 0.010587, 0.010582, 0.010577, 
    0.010572, 0.010567, 0.010563, 0.010558, 0.010553, 0.010547, 0.010542, 
    0.010536, 0.01053, 0.010524, 0.010518, 0.010512, 0.010505, 0.010497, 
    0.010488, 0.010479, 0.01047, 0.010464, 0.010458, 0.010452, 0.010446, 
    0.010439, 0.010431, 0.010423, 0.010412, 0.010402, 0.010394, 0.010387, 
    0.01038, 0.010369, 0.010358, 0.010345, 0.010333, 0.010321, 0.010311, 
    0.010301, 0.010292, 0.010283, 0.010274, 0.010266, 0.010259, 0.010252, 
    0.010245, 0.010238, 0.010231, 0.010224, 0.010218, 0.01021, 0.010202, 
    0.010196, 0.010189, 0.010183, 0.010178, 0.010174, 0.010169, 0.010162, 
    0.010156, 0.010148, 0.010141, 0.010134, 0.010128, 0.010124, 0.01012, 
    0.010115, 0.010111, 0.010108, 0.010103, 0.010102, 0.010103, 0.010105, 
    0.010107, 0.01011, 0.010112, 0.010112, 0.010113, 0.010113, 0.010114, 
    0.010114, 0.010115, 0.010117, 0.010119, 0.01012, 0.010121, 0.010122, 
    0.010123, 0.010123, 0.010124, 0.010126, 0.010128, 0.010129, 0.010131, 
    0.010132, 0.010132, 0.010134, 0.010136, 0.010139, 0.010142, 0.010146, 
    0.010149, 0.010151, 0.010154, 0.010156, 0.010158, 0.010159, 0.01016, 
    0.010163, 0.010163, 0.010162, 0.010159, 0.010156, 0.010153, 0.010152, 
    0.010152, 0.010152, 0.010151, 0.01015, 0.010149, 0.010148, 0.010147, 
    0.010146, 0.010145, 0.010144, 0.010143, 0.010144, 0.010144, 0.010143, 
    0.010143, 0.010143, 0.010142, 0.010142, 0.010143, 0.010143, 0.010141, 
    0.01014, 0.010138, 0.010135, 0.010133, 0.010131, 0.010129, 0.010126, 
    0.010123, 0.01012, 0.010115, 0.01011, 0.010106, 0.010105, 0.010104, 
    0.010105, 0.010106, 0.010106, 0.010103, 0.010099, 0.010097, 0.010095, 
    0.010093, 0.010092, 0.010089, 0.010086, 0.010079, 0.010072, 0.010065, 
    0.010058, 0.010052, 0.010048, 0.010045, 0.010042, 0.010039, 0.010035, 
    0.010031, 0.010026, 0.010021, 0.010016, 0.010013, 0.010012, 0.010011, 
    0.010006, 0.01, 0.0099963, 0.0099919, 0.0099869, 0.0099846, 0.0099827, 
    0.0099798, 0.0099758, 0.0099705, 0.0099629, 0.0099545, 0.0099459, 
    0.0099387, 0.0099337, 0.0099277, 0.0099214, 0.0099155, 0.0099089, 
    0.0099006, 0.009894, 0.0098882, 0.0098872, 0.0098861, 0.0098846, 
    0.0098834, 0.0098824, 0.0098783, 0.0098739, 0.0098688, 0.0098633, 
    0.0098574, 0.0098547, 0.0098527, 0.0098521, 0.009849, 0.0098436, 
    0.009837, 0.0098304, 0.0098248, 0.0098198, 0.0098153, 0.0098113, 
    0.0098076, 0.0098038, 0.0097988, 0.0097921, 0.0097864, 0.0097813, 
    0.00978, 0.0097788, 0.0097776, 0.0097766, 0.0097756, 0.0097727, 
    0.0097701, 0.0097679, 0.0097669, 0.0097665, 0.0097674, 0.0097675, 
    0.0097657, 0.009763, 0.0097598, 0.0097534, 0.0097467, 0.0097396, 
    0.0097363, 0.009736, 0.0097321, 0.009727, 0.0097189, 0.0097102, 
    0.0097011, 0.0096947, 0.0096893, 0.0096859, 0.0096822, 0.0096781, 
    0.0096742, 0.00967, 0.0096644, 0.009659, 0.0096539, 0.0096525, 0.0096521, 
    0.0096508, 0.0096488, 0.0096458, 0.00964, 0.0096332, 0.0096273, 
    0.0096211, 0.0096144, 0.0096076, 0.0096007, 0.0095942, 0.0095878, 
    0.0095816, 0.0095759, 0.0095706, 0.0095653, 0.0095602, 0.009556, 
    0.0095524, 0.0095493, 0.0095417, 0.0095347, 0.0095329, 0.0095306, 
    0.0095278, 0.0095246, 0.0095215, 0.0095184, 0.0095154, 0.0095127, 
    0.0095107, 0.0095088, 0.0095059, 0.0095033, 0.0095012, 0.0094965, 
    0.0094908, 0.009484, 0.0094772, 0.0094703, 0.0094656, 0.009462, 
    0.0094606, 0.0094592, 0.0094578, 0.0094574, 0.0094576, 0.009456, 
    0.0094541, 0.0094516, 0.0094481, 0.0094441, 0.0094404, 0.0094366, 
    0.0094325, 0.009429, 0.0094259, 0.0094219, 0.0094175, 0.0094123, 
    0.0094079, 0.0094042, 0.0094017, 0.0093994, 0.0093972, 0.0093944, 
    0.0093909, 0.0093874, 0.0093841, 0.0093815, 0.0093799, 0.0093796, 
    0.0093789, 0.0093782, 0.0093791, 0.0093801, 0.0093815, 0.0093819, 
    0.0093819, 0.0093812, 0.0093799, 0.0093775, 0.0093739, 0.0093698, 
    0.0093656, 0.0093615, 0.0093578, 0.0093527, 0.0093467, 0.0093403, 
    0.0093343, 0.0093298, 0.0093257, 0.0093221, 0.0093185, 0.009315, 
    0.0093123, 0.0093093, 0.0093062, 0.0093021, 0.0092979, 0.0092943, 
    0.0092905, 0.0092864, 0.0092833, 0.0092804, 0.0092772, 0.0092734, 
    0.0092686, 0.009264, 0.0092596, 0.0092562, 0.0092524, 0.0092477, 
    0.0092427, 0.0092376, 0.0092324, 0.0092273, 0.0092222, 0.0092162, 
    0.0092097, 0.0092028, 0.0091952, 0.0091862, 0.0091781, 0.0091705, 
    0.009168, 0.0091661, 0.0091646, 0.0091628, 0.0091607, 0.0091575, 
    0.0091538, 0.0091491, 0.0091446, 0.0091405, 0.0091362, 0.0091322, 
    0.0091301, 0.0091275, 0.0091243, 0.0091215, 0.0091186, 0.0091145, 
    0.0091105, 0.0091067, 0.0091025, 0.0090982, 0.0090927, 0.0090876, 
    0.009083, 0.0090776, 0.0090719, 0.0090657, 0.0090595, 0.0090533, 
    0.0090474, 0.0090417, 0.0090383, 0.0090359, 0.0090353, 0.0090354, 
    0.009036, 0.009035, 0.0090335, 0.0090304, 0.0090273, 0.0090242, 
    0.0090207, 0.0090176, 0.0090159, 0.009014, 0.0090118, 0.009008, 
    0.0090035, 0.0089968, 0.0089898, 0.0089826, 0.0089771, 0.0089723, 
    0.0089701, 0.0089678, 0.0089655, 0.0089606, 0.008955, 0.0089515, 
    0.0089486, 0.0089468, 0.0089483, 0.0089512, 0.0089507, 0.00895, 
    0.0089493, 0.008948, 0.0089463, 0.0089453, 0.0089443, 0.008943, 
    0.0089415, 0.0089397, 0.0089388, 0.008938, 0.0089369, 0.0089359, 
    0.0089349, 0.0089331, 0.0089313, 0.0089297, 0.0089276, 0.0089249, 
    0.0089239, 0.0089235, 0.0089245, 0.0089262, 0.0089284, 0.0089305, 
    0.0089322, 0.0089315, 0.0089296, 0.0089261, 0.0089227, 0.0089196, 
    0.0089212, 0.00892, 0.0089147, 0.0089075, 0.0088994, 0.0088896, 
    0.0088812, 0.0088753, 0.0088701, 0.0088652, 0.008862, 0.0088585, 
    0.0088538, 0.0088487, 0.0088435, 0.008841, 0.0088388, 0.0088368, 
    0.008834, 0.0088305, 0.0088254, 0.00882, 0.0088145, 0.0088093, 0.0088044, 
    0.0088017, 0.0087993, 0.0087953, 0.0087915, 0.008788, 0.008784, 
    0.0087798, 0.0087752, 0.0087709, 0.0087671, 0.0087646, 0.0087623, 
    0.008759, 0.0087557, 0.0087525, 0.0087506, 0.0087492, 0.0087492, 
    0.0087489, 0.0087482, 0.008748, 0.0087482, 0.0087483, 0.008749, 
    0.0087514, 0.0087545, 0.0087581, 0.00876, 0.0087614, 0.008762, 0.0087614, 
    0.0087599, 0.00876, 0.0087606, 0.0087623, 0.0087629, 0.0087627, 
    0.0087614, 0.0087597, 0.0087564, 0.0087541, 0.0087527, 0.0087512, 
    0.0087498, 0.0087488, 0.0087482, 0.008748, 0.0087465, 0.0087445, 
    0.0087428, 0.0087411, 0.0087394, 0.0087385, 0.0087379, 0.0087375, 
    0.0087365, 0.0087342, 0.0087329, 0.008732, 0.0087308, 0.0087291, 
    0.0087264, 0.0087227, 0.0087186, 0.0087137, 0.0087088, 0.0087038, 
    0.0086995, 0.0086958, 0.0086928, 0.0086897, 0.0086852, 0.0086804, 
    0.0086754, 0.0086703, 0.0086653, 0.0086603, 0.0086552, 0.0086499, 
    0.0086442, 0.0086383, 0.0086323, 0.0086263, 0.0086202, 0.0086146, 
    0.0086095, 0.0086069, 0.0086043, 0.0086018, 0.008599, 0.008596, 0.008594, 
    0.0085923, 0.0085913, 0.0085892, 0.0085865, 0.0085819, 0.0085774, 
    0.0085735, 0.0085688, 0.0085636, 0.0085606, 0.0085581, 0.0085568, 
    0.0085554, 0.0085541, 0.0085489, 0.0085432, 0.008537, 0.0085318, 
    0.0085275, 0.0085236, 0.0085201, 0.0085182, 0.0085166, 0.0085154, 
    0.0085143, 0.0085133, 0.0085132, 0.0085132, 0.0085134, 0.0085125, 
    0.0085111, 0.0085086, 0.0085051, 0.0084998, 0.0084966, 0.0084942, 
    0.008491, 0.0084868, 0.0084808, 0.0084757, 0.0084711, 0.0084705, 
    0.0084707, 0.0084727, 0.0084734, 0.0084733, 0.0084743, 0.0084745, 
    0.0084724, 0.0084699, 0.008467, 0.0084647, 0.0084627, 0.0084621, 
    0.0084621, 0.0084626, 0.0084638, 0.0084653, 0.0084672, 0.008469, 
    0.0084707, 0.0084715, 0.0084719, 0.0084719, 0.0084709, 0.0084685, 
    0.0084671, 0.008466, 0.0084638, 0.0084611, 0.0084576, 0.0084536, 
    0.0084495, 0.0084462, 0.0084433, 0.0084412, 0.0084401, 0.0084394, 
    0.0084389, 0.0084376, 0.0084342, 0.0084308, 0.0084275, 0.0084242, 
    0.0084209, 0.0084179, 0.0084148, 0.0084117, 0.0084089, 0.0084058, 
    0.0084014, 0.0083974, 0.0083939, 0.0083888, 0.0083832, 0.0083766, 
    0.0083695, 0.0083619, 0.0083545, 0.0083472, 0.0083403, 0.0083339, 
    0.0083282, 0.0083232, 0.0083184, 0.0083128, 0.0083083, 0.0083054, 
    0.0083041, 0.0083034, 0.0083021, 0.0082999, 0.0082963, 0.0082925, 
    0.0082887, 0.0082838, 0.008278, 0.0082701, 0.008262, 0.0082538, 
    0.0082455, 0.0082372, 0.0082291, 0.0082211, 0.0082132, 0.0082052, 
    0.008197, 0.0081882, 0.0081811, 0.0081755, 0.008171, 0.0081671, 
    0.0081656, 0.0081636, 0.0081612, 0.0081591, 0.008157, 0.0081552, 
    0.0081535, 0.0081518, 0.0081499, 0.0081479, 0.0081446, 0.0081413, 
    0.008138, 0.0081335, 0.0081285, 0.0081234, 0.0081185, 0.0081137, 
    0.0081092, 0.0081049, 0.0081019, 0.0080992, 0.0080974, 0.008097, 
    0.0080975, 0.0080982, 0.008099, 0.0081001, 0.0081006, 0.0081006, 
    0.0080987, 0.0080969, 0.0080962, 0.0080955, 0.0080949, 0.0080926, 
    0.0080898, 0.0080861, 0.0080816, 0.0080762, 0.0080717, 0.0080675, 
    0.0080646, 0.0080624, 0.0080609, 0.0080595, 0.008058, 0.008057, 
    0.0080563, 0.0080561, 0.0080562, 0.0080564, 0.0080572, 0.0080572, 
    0.0080559, 0.0080557, 0.008056, 0.0080547, 0.0080532, 0.0080513, 
    0.0080495, 0.008048, 0.0080476, 0.0080471, 0.0080462, 0.0080455, 
    0.0080449, 0.0080454, 0.0080461, 0.008047, 0.0080478, 0.0080484, 
    0.0080478, 0.008047, 0.0080462, 0.0080449, 0.0080432, 0.0080427, 
    0.0080428, 0.0080445, 0.0080459, 0.0080468, 0.0080471, 0.008047, 
    0.0080456, 0.0080447, 0.0080444, 0.0080435, 0.0080424, 0.0080414, 
    0.0080397, 0.0080368, 0.0080344, 0.0080321, 0.0080312, 0.0080311, 
    0.0080328, 0.0080334, 0.0080334, 0.0080321, 0.0080304, 0.008028, 
    0.0080259, 0.0080239, 0.0080217, 0.0080193, 0.0080168, 0.0080142, 
    0.0080116, 0.008009, 0.0080069, 0.0080075, 0.0080084, 0.0080096, 
    0.0080107, 0.0080117, 0.0080125, 0.0080123, 0.008011, 0.00801, 0.008009, 
    0.0080071, 0.0080048, 0.0080021, 0.0079993, 0.0079967, 0.007994, 
    0.0079916, 0.0079895, 0.0079886, 0.0079883, 0.0079867, 0.0079844, 
    0.0079805, 0.0079759, 0.0079708, 0.0079666, 0.0079625, 0.007958, 
    0.0079536, 0.0079491, 0.0079443, 0.0079397, 0.0079357, 0.0079325, 
    0.0079301, 0.0079275, 0.0079248, 0.0079214, 0.0079177, 0.0079138, 
    0.0079102, 0.007907, 0.0079059, 0.0079045, 0.0079026, 0.0078997, 
    0.0078964, 0.0078918, 0.007888, 0.0078857, 0.0078845, 0.0078836, 
    0.0078815, 0.0078798, 0.0078787, 0.0078774, 0.0078761, 0.0078742, 
    0.0078724, 0.0078708, 0.0078692, 0.0078676, 0.0078669, 0.0078662, 
    0.0078653, 0.0078644, 0.0078634, 0.0078618, 0.0078604, 0.0078596, 
    0.0078586, 0.0078574, 0.0078556, 0.0078536, 0.0078509, 0.0078478, 
    0.0078444, 0.0078417, 0.0078392, 0.007837, 0.0078341, 0.0078303, 
    0.0078269, 0.0078238, 0.0078209, 0.0078182, 0.0078156, 0.0078132, 
    0.007811, 0.0078086, 0.0078063, 0.0078043, 0.0078021, 0.0077996, 
    0.0077968, 0.0077942, 0.0077923, 0.0077904, 0.0077885, 0.0077868, 
    0.0077846, 0.007781, 0.0077777, 0.0077747, 0.0077721, 0.0077693, 
    0.0077659, 0.0077625, 0.0077592, 0.0077561, 0.0077533, 0.0077514, 
    0.0077498, 0.0077487, 0.0077475, 0.0077459, 0.007742, 0.0077379, 
    0.0077337, 0.0077305, 0.0077275, 0.0077234, 0.007719, 0.0077139, 
    0.0077086, 0.0077032, 0.0076974, 0.0076916, 0.0076858, 0.0076793, 
    0.0076725, 0.007667, 0.0076617, 0.0076567, 0.0076522, 0.007648, 
    0.0076442, 0.0076408, 0.0076381, 0.0076363, 0.0076352, 0.007635, 
    0.0076349, 0.0076349, 0.0076341, 0.0076327, 0.0076297, 0.0076263, 
    0.0076218, 0.0076177, 0.0076141, 0.0076108, 0.0076075, 0.0076031, 
    0.007599, 0.0075951, 0.0075903, 0.0075853, 0.007581, 0.0075777, 
    0.0075758, 0.007574, 0.0075722, 0.0075704, 0.0075683, 0.007566, 
    0.0075645, 0.0075633, 0.0075631, 0.007563, 0.0075631, 0.0075628, 
    0.0075623, 0.0075602, 0.0075579, 0.007555, 0.0075518, 0.0075483, 
    0.0075454, 0.007542, 0.007537, 0.0075322, 0.0075275, 0.0075253, 
    0.0075239, 0.0075234, 0.0075232, 0.0075233, 0.007522, 0.0075205, 
    0.0075195, 0.0075182, 0.0075165, 0.0075169, 0.0075177, 0.0075152, 
    0.0075123, 0.0075087, 0.0075065, 0.0075049, 0.0075025, 0.0075008, 
    0.0075001, 0.0075011, 0.0075029, 0.0075045, 0.0075055, 0.0075052, 
    0.0075046, 0.0075038, 0.0075022, 0.0075006, 0.0074994, 0.0074981, 
    0.0074967, 0.0074942, 0.0074912, 0.0074865, 0.0074831, 0.0074809, 
    0.0074797, 0.0074784, 0.0074758, 0.0074732, 0.0074704, 0.0074679, 
    0.0074655, 0.007464, 0.0074626, 0.0074615, 0.0074614, 0.0074615, 
    0.0074607, 0.0074609, 0.0074624, 0.0074637, 0.0074648, 0.0074635, 
    0.0074629, 0.0074635, 0.0074618, 0.0074589, 0.0074538, 0.0074486, 
    0.0074434, 0.0074382, 0.0074329, 0.0074286, 0.0074247, 0.0074217, 
    0.0074187, 0.0074158, 0.0074134, 0.0074111, 0.0074092, 0.0074076, 
    0.0074062, 0.0074042, 0.0074017, 0.0073982, 0.0073964, 0.0073965, 
    0.0073979, 0.0073994, 0.0073987, 0.0073966, 0.0073927, 0.0073896, 
    0.0073869, 0.0073843, 0.0073821, 0.0073806, 0.0073788, 0.007377, 
    0.007374, 0.0073713, 0.0073692, 0.0073676, 0.0073662, 0.007366, 
    0.0073657, 0.0073648, 0.0073639, 0.0073631, 0.0073633, 0.0073637, 
    0.007364, 0.0073648, 0.0073659, 0.0073663, 0.0073664, 0.0073653, 
    0.0073641, 0.0073626, 0.0073615, 0.0073604, 0.0073596, 0.0073589, 
    0.0073582, 0.0073542, 0.0073493, 0.0073438, 0.0073396, 0.0073371, 
    0.0073361, 0.0073356, 0.0073352, 0.0073344, 0.0073327, 0.0073299, 
    0.0073266, 0.0073225, 0.0073188, 0.0073159, 0.0073127, 0.0073092, 
    0.0073051, 0.0073012, 0.0072982, 0.0072954, 0.0072929, 0.0072914, 
    0.0072898, 0.007288, 0.0072862, 0.0072845, 0.0072828, 0.0072815, 
    0.0072818, 0.0072824, 0.0072831, 0.0072835, 0.0072838, 0.0072838, 
    0.0072839, 0.007284, 0.007284, 0.0072841, 0.0072846, 0.0072853, 0.007286, 
    0.0072867, 0.0072873, 0.0072883, 0.0072898, 0.0072918, 0.0072942, 
    0.0072969, 0.0073012, 0.0073057, 0.0073108, 0.0073156, 0.0073204, 
    0.0073248, 0.0073286, 0.007331, 0.0073326, 0.0073337, 0.0073345, 
    0.0073352, 0.0073357, 0.0073364, 0.0073372, 0.0073393, 0.0073412, 
    0.0073422, 0.0073428, 0.0073431, 0.0073451, 0.0073474, 0.0073498, 
    0.0073522, 0.0073546, 0.007357, 0.0073594, 0.007362, 0.0073642, 
    0.0073657, 0.0073677, 0.0073698, 0.0073714, 0.0073729, 0.0073743, 
    0.0073753, 0.0073761, 0.007376, 0.0073752, 0.0073733, 0.0073712, 
    0.0073691, 0.0073679, 0.0073669, 0.0073663, 0.0073671, 0.0073687, 
    0.0073693, 0.0073694, 0.0073687, 0.0073682, 0.007368, 0.0073671, 
    0.007366, 0.0073646, 0.0073643, 0.0073651, 0.0073662, 0.0073671, 
    0.0073673, 0.0073675, 0.0073678, 0.0073674, 0.0073667, 0.0073647, 
    0.0073625, 0.0073599, 0.0073571, 0.0073543, 0.0073509, 0.0073471, 
    0.0073428, 0.0073384, 0.007334, 0.0073302, 0.0073272, 0.0073259, 
    0.0073257, 0.0073261, 0.0073262, 0.0073259, 0.0073246, 0.0073229, 
    0.0073211, 0.0073195, 0.0073181, 0.0073172, 0.0073166, 0.0073161, 
    0.0073144, 0.0073125, 0.0073103, 0.0073072, 0.0073035, 0.0072983, 
    0.0072928, 0.0072873, 0.0072818, 0.0072764, 0.0072715, 0.007267, 
    0.007264, 0.0072617, 0.0072603, 0.00726, 0.0072602, 0.0072612, 0.0072624, 
    0.0072636, 0.0072645, 0.0072652, 0.0072647, 0.007264, 0.0072627, 
    0.0072598, 0.0072562, 0.0072523, 0.0072485, 0.0072448, 0.0072415, 
    0.0072386, 0.0072361, 0.0072335, 0.0072306, 0.0072281, 0.007226, 
    0.0072238, 0.0072215, 0.0072187, 0.007216, 0.0072133, 0.0072105, 
    0.0072079, 0.0072058, 0.007203, 0.0071994, 0.0071959, 0.0071923, 
    0.0071883, 0.007184, 0.007179, 0.0071741, 0.007169, 0.0071634, 0.0071583, 
    0.0071539, 0.0071483, 0.0071422, 0.0071382, 0.0071341, 0.0071296, 
    0.0071247, 0.0071196, 0.0071145, 0.007109, 0.0071025, 0.0070954, 
    0.0070879, 0.0070805, 0.0070733, 0.0070664, 0.0070596, 0.0070527, 
    0.0070474, 0.0070425, 0.0070385, 0.0070348, 0.0070315, 0.0070284, 
    0.0070252, 0.0070216, 0.0070167, 0.0070103, 0.0070051, 0.0069999, 
    0.006994, 0.0069875, 0.0069804, 0.0069719, 0.0069628, 0.0069523, 
    0.0069416, 0.0069303, 0.0069189, 0.0069073, 0.0068951, 0.0068821, 
    0.0068674, 0.006853, 0.0068387, 0.0068246, 0.0068109, 0.006798, 
    0.0067868, 0.0067767, 0.0067659, 0.0067551, 0.0067442, 0.006733, 
    0.0067217, 0.0067103, 0.0066988, 0.0066869, 0.0066744, 0.0066613, 
    0.0066483, 0.0066354, 0.0066228, 0.0066111, 0.0066002, 0.0065915, 
    0.0065834, 0.0065755, 0.0065678, 0.0065604, 0.006555, 0.0065503, 
    0.0065468, 0.0065426, 0.0065372, 0.0065324, 0.0065279, 0.006525, 
    0.0065228, 0.0065218, 0.0065216, 0.0065218, 0.0065222, 0.0065224, 
    0.0065223, 0.0065223, 0.0065223, 0.0065228, 0.0065236, 0.0065249, 
    0.0065257, 0.0065262, 0.0065275, 0.0065288, 0.00653, 0.0065306, 
    0.0065308, 0.0065317, 0.0065324, 0.006531, 0.0065292, 0.0065268, 
    0.0065243, 0.0065216, 0.0065176, 0.0065134, 0.0065089, 0.006505, 
    0.0065012, 0.006497, 0.0064936, 0.0064911, 0.0064914, 0.0064927, 
    0.0064923, 0.0064915, 0.0064901, 0.006489, 0.006488, 0.0064869, 
    0.0064865, 0.0064875, 0.0064891, 0.006491, 0.0064907, 0.0064898, 
    0.0064872, 0.0064852, 0.0064835, 0.0064836, 0.006484, 0.0064852, 
    0.0064854, 0.0064848, 0.0064841, 0.0064838, 0.006485, 0.0064873, 
    0.0064908, 0.0064944, 0.0064982, 0.0065021, 0.0065062, 0.0065104, 
    0.0065146, 0.006519, 0.0065238, 0.0065286, 0.0065334, 0.0065377, 
    0.0065418, 0.0065458, 0.00655, 0.0065548, 0.0065591, 0.0065631, 
    0.0065679, 0.0065724, 0.0065763, 0.0065793, 0.0065817, 0.0065832, 
    0.0065845, 0.0065856, 0.0065873, 0.0065895, 0.0065896, 0.0065885, 
    0.0065841, 0.0065794, 0.0065744, 0.0065708, 0.0065673, 0.0065633, 
    0.0065589, 0.0065541, 0.0065501, 0.0065463, 0.0065425, 0.0065388, 
    0.0065353, 0.006532, 0.0065287, 0.0065245, 0.0065205, 0.0065165, 
    0.0065127, 0.0065091, 0.006504, 0.0064985, 0.0064921, 0.0064857, 
    0.0064791, 0.0064732, 0.0064675, 0.006462, 0.0064574, 0.0064533, 
    0.0064482, 0.0064433, 0.0064386, 0.0064348, 0.0064316, 0.006429, 
    0.0064266, 0.0064244, 0.0064229, 0.0064221, 0.0064214, 0.0064207, 
    0.0064201, 0.0064196, 0.0064193, 0.0064198, 0.0064204, 0.0064201, 
    0.0064195, 0.0064187, 0.0064178, 0.0064169, 0.0064161, 0.0064145, 
    0.0064117, 0.0064068, 0.0064009, 0.0063933, 0.0063857, 0.0063779, 
    0.0063699, 0.0063619, 0.0063537, 0.0063453, 0.0063363, 0.0063269, 
    0.0063172, 0.0063084, 0.0063003, 0.0062936, 0.0062883, 0.0062842, 
    0.0062803, 0.0062765, 0.0062725, 0.0062678, 0.0062626, 0.0062571, 
    0.0062516, 0.0062461, 0.0062405, 0.0062348, 0.0062287, 0.0062224, 
    0.0062147, 0.0062075, 0.0062006, 0.0061944, 0.0061885, 0.0061839, 
    0.0061803, 0.0061782, 0.0061781, 0.0061788, 0.0061813, 0.0061844, 
    0.0061884, 0.0061931, 0.0061981, 0.0062027, 0.0062065, 0.0062088, 
    0.0062101, 0.0062108, 0.0062111, 0.006211, 0.0062099, 0.006208, 
    0.0062053, 0.0062013, 0.0061969, 0.0061919, 0.0061865, 0.0061809, 
    0.0061775, 0.0061744, 0.0061713, 0.0061677, 0.0061637, 0.0061595, 
    0.0061552, 0.0061504, 0.0061457, 0.006141, 0.0061365, 0.0061319, 
    0.0061259, 0.006119, 0.0061106, 0.0061016, 0.0060922, 0.0060839, 
    0.0060759, 0.0060684, 0.0060615, 0.0060549, 0.0060492, 0.0060439, 
    0.0060395, 0.0060359, 0.0060329, 0.0060302, 0.0060276, 0.0060249, 
    0.0060213, 0.006017, 0.0060123, 0.0060075, 0.0060033, 0.0059991, 
    0.0059949, 0.0059913, 0.0059878, 0.0059843, 0.0059805, 0.0059766, 
    0.0059734, 0.0059704, 0.0059674, 0.0059647, 0.0059622, 0.0059586, 
    0.0059545, 0.0059501, 0.0059457, 0.0059412, 0.0059367, 0.0059322, 
    0.0059278, 0.0059225, 0.0059154, 0.0059073, 0.0058988, 0.0058886, 
    0.0058778, 0.0058657, 0.0058537, 0.0058416, 0.0058314, 0.0058219, 
    0.0058141, 0.005807, 0.0058004, 0.0057959, 0.0057917, 0.0057878, 
    0.0057839, 0.0057801, 0.0057767, 0.0057734, 0.0057695, 0.0057652, 
    0.0057605, 0.0057558, 0.0057511, 0.0057459, 0.0057404, 0.0057347, 
    0.0057289, 0.0057232, 0.005718, 0.0057129, 0.005708, 0.005703, 0.0056978, 
    0.0056919, 0.0056855, 0.0056779, 0.0056707, 0.0056636, 0.0056572, 
    0.005651, 0.0056456, 0.0056404, 0.0056354, 0.0056298, 0.0056241, 
    0.005618, 0.0056114, 0.0056042, 0.0055982, 0.0055922, 0.0055857, 
    0.0055792, 0.0055726, 0.0055658, 0.0055589, 0.0055522, 0.0055458, 
    0.0055397, 0.0055341, 0.0055287, 0.0055237, 0.0055188, 0.0055142, 
    0.0055094, 0.0055044, 0.0054991, 0.0054939, 0.0054889, 0.0054851, 
    0.0054819, 0.0054803, 0.0054793, 0.0054796, 0.0054801, 0.0054806, 
    0.0054825, 0.0054845, 0.0054866, 0.0054891, 0.0054919, 0.0054959, 
    0.0054999, 0.0055038, 0.0055067, 0.0055088, 0.0055098, 0.0055107, 
    0.005512, 0.0055133, 0.0055147, 0.0055159, 0.0055168, 0.0055162, 
    0.0055142, 0.0055107, 0.005507, 0.0055032, 0.0054994, 0.0054956, 
    0.0054918, 0.0054882, 0.0054847, 0.0054824, 0.0054804, 0.0054791, 
    0.005478, 0.0054769, 0.0054747, 0.0054724, 0.0054697, 0.005467, 
    0.0054643, 0.0054618, 0.0054591, 0.005456, 0.0054523, 0.0054484, 
    0.0054432, 0.0054375, 0.0054308, 0.0054247, 0.005419, 0.0054148, 
    0.0054105, 0.0054056, 0.0054003, 0.0053945, 0.0053882, 0.0053818, 
    0.0053755, 0.0053704, 0.0053667, 0.0053649, 0.0053636, 0.0053622, 
    0.0053605, 0.0053587, 0.0053567, 0.0053548, 0.0053527, 0.0053505, 
    0.0053482, 0.0053455, 0.0053426, 0.0053387, 0.0053345, 0.00533, 
    0.0053251, 0.00532, 0.0053142, 0.005308, 0.0053012, 0.0052939, 0.0052863, 
    0.0052796, 0.0052731, 0.0052668, 0.0052607, 0.0052548, 0.0052487, 
    0.0052425, 0.0052359, 0.0052292, 0.0052224, 0.0052152, 0.0052081, 
    0.0052017, 0.0051952, 0.0051887, 0.0051816, 0.0051744, 0.0051674, 
    0.0051608, 0.0051549, 0.0051501, 0.0051459, 0.0051427, 0.0051398, 
    0.0051373, 0.0051347, 0.0051323, 0.0051302, 0.0051282, 0.0051266, 
    0.0051249, 0.0051231, 0.0051213, 0.0051195, 0.005118, 0.0051161, 
    0.0051139, 0.0051121, 0.00511, 0.0051073, 0.0051047, 0.0051021, 
    0.0050995, 0.0050969, 0.0050946, 0.0050925, 0.0050906, 0.0050891, 
    0.0050877, 0.0050865, 0.0050852, 0.005084, 0.0050833, 0.0050828, 
    0.0050824, 0.005082, 0.0050815, 0.0050809, 0.0050801, 0.0050773, 
    0.0050741, 0.0050702, 0.0050665, 0.0050628, 0.0050582, 0.0050533, 
    0.0050478, 0.0050424, 0.0050373, 0.0050319, 0.0050267, 0.0050221, 
    0.0050183, 0.0050152, 0.0050129, 0.0050107, 0.0050083, 0.0050063, 
    0.0050045, 0.0050022, 0.0049996, 0.0049959, 0.0049919, 0.0049878, 
    0.0049831, 0.0049781, 0.0049722, 0.0049664, 0.0049607, 0.0049552, 
    0.0049498, 0.0049442, 0.0049389, 0.0049337, 0.0049284, 0.004923, 
    0.0049175, 0.0049123, 0.0049074, 0.0049029, 0.0048984, 0.0048939, 
    0.0048892, 0.0048839, 0.0048784, 0.0048728, 0.0048673, 0.0048624, 
    0.0048585, 0.0048544, 0.0048502, 0.004845, 0.0048398, 0.0048348, 
    0.0048295, 0.004824, 0.0048191, 0.0048144, 0.0048104, 0.0048071, 
    0.0048043, 0.0048016, 0.004799, 0.0047967, 0.0047948, 0.0047933, 
    0.0047921, 0.004791, 0.00479, 0.004789, 0.0047879, 0.0047859, 0.0047836, 
    0.0047809, 0.0047779, 0.0047745, 0.0047711, 0.0047677, 0.0047639, 
    0.0047602, 0.004757, 0.0047547, 0.0047529, 0.0047511, 0.0047493, 
    0.0047759, 0.004766, 0.0047561, 0.0047461, 0.0047361, 0.004726, 
    0.0047159, 0.0047058, 0.0046957, 0.0046856, 0.0046755, 0.0046654, 
    0.0046553, 0.0046454, 0.0046355, 0.0046256, 0.0046159, 0.0046062, 
    0.0045967, 0.0045873, 0.004578, 0.0045688, 0.0045597, 0.0045507, 
    0.0045418, 0.0045331, 0.0045244, 0.0045157, 0.0045072, 0.0044987, 
    0.0044902, 0.0044817, 0.0044732, 0.0044648, 0.0044563, 0.0044478, 
    0.0044392, 0.0044306, 0.004422, 0.0044133, 0.0044046, 0.0043959, 
    0.0043871, 0.0043783, 0.0043694, 0.0043606, 0.0043517, 0.0043428, 
    0.004334, 0.0043251, 0.0043163, 0.0043075, 0.0042987, 0.0042899, 
    0.0042812, 0.0042725, 0.0042639, 0.0042553, 0.0042467, 0.0042382, 
    0.0042297, 0.0042212, 0.0042127, 0.0042042, 0.0041957, 0.0041872, 
    0.0041787, 0.0041701, 0.0041615, 0.0041529, 0.0041442, 0.0041355, 
    0.0041267, 0.0041179, 0.004109, 0.0041001, 0.0040911, 0.0040821, 
    0.004073, 0.0040639, 0.0040548, 0.0040456, 0.0040364, 0.0040272, 
    0.004018, 0.0040088, 0.0039995, 0.0039903, 0.0039811, 0.0039719, 
    0.0039627, 0.0039535, 0.0039443, 0.0039352, 0.003926, 0.0039169, 
    0.0039078, 0.0038987, 0.0038896, 0.0038805, 0.0038714, 0.0038623, 
    0.0038532, 0.0038441, 0.0038351, 0.003826, 0.003817, 0.0038079, 
    0.0037988, 0.0037898, 0.0037807, 0.0037717, 0.0037626, 0.0037536, 
    0.0037445, 0.0037355, 0.0037264, 0.0037174, 0.0037083, 0.0036992, 
    0.0036902, 0.0036811, 0.003672, 0.003663, 0.0036539, 0.0036448, 
    0.0036357, 0.0036266, 0.0036175, 0.0036084, 0.0035993, 0.0035902, 
    0.0035811, 0.003572, 0.003563, 0.0035539, 0.0035448, 0.0035358, 
    0.0035267, 0.0035177, 0.0035087, 0.0034997, 0.0034908, 0.0034819, 
    0.003473, 0.0034642, 0.0034554, 0.0034467, 0.003438, 0.0034294, 
    0.0034208, 0.0034123, 0.0034039, 0.0033955, 0.0033871, 0.0033789, 
    0.0033706, 0.0033625, 0.0033543, 0.0033462, 0.0033382, 0.0033302, 
    0.0033222, 0.0033143, 0.0033064, 0.0032985, 0.0032907, 0.0032828, 
    0.003275, 0.0032672, 0.0032594, 0.0032517, 0.0032439, 0.0032361, 
    0.0032284, 0.0032206, 0.0032129, 0.0032051, 0.0031974, 0.0031896, 
    0.0031819, 0.0031741, 0.0031664, 0.0031586, 0.0031509, 0.0031431, 
    0.0031354, 0.0031276, 0.0031199, 0.0031121, 0.0031044, 0.0030966, 
    0.0030888, 0.0030811, 0.0030733, 0.0030655, 0.0030577, 0.0030499, 
    0.0030421, 0.0030343, 0.0030266, 0.0030188, 0.003011, 0.0030033, 
    0.0029956, 0.0029879, 0.0029802, 0.0029726, 0.0029651, 0.0029576, 
    0.0029502, 0.0029428, 0.0029355, 0.0029283, 0.0029211, 0.0029141, 
    0.0029071, 0.0029001, 0.0028933, 0.0028865, 0.0028797, 0.002873, 
    0.0028663, 0.0028597, 0.0028531, 0.0028465, 0.00284, 0.0028334, 
    0.0028269, 0.0028204, 0.0028138, 0.0028072, 0.0028006, 0.002794, 
    0.0027874, 0.0027808, 0.0027741, 0.0027674, 0.0027607, 0.002754, 
    0.0027472, 0.0027404, 0.0027337, 0.0027269, 0.00272, 0.0027132, 
    0.0027063, 0.0026994, 0.0026925, 0.0026856, 0.0026786, 0.0026716, 
    0.0026646, 0.0026575, 0.0026504, 0.0026432, 0.002636, 0.0026287, 
    0.0026214, 0.002614, 0.0026066, 0.002599, 0.0025915, 0.0025838, 
    0.0025761, 0.0025684, 0.0025606, 0.0025527, 0.0025448, 0.0025368, 
    0.0025288, 0.0025208, 0.0025128, 0.0025048, 0.0024967, 0.0024887, 
    0.0024807, 0.0024726, 0.0024647, 0.0024567, 0.0024488, 0.002441, 
    0.0024332, 0.0024254, 0.0024177, 0.00241, 0.0024024, 0.0023948, 
    0.0023873, 0.0023798, 0.0023723, 0.0023648, 0.0023574, 0.00235, 
    0.0023427, 0.0023353, 0.002328, 0.0023207, 0.0023134, 0.0023062, 
    0.0022989, 0.0022918, 0.0022846, 0.0022776, 0.0022706, 0.0022636, 
    0.0022567, 0.0022499, 0.0022431, 0.0022364, 0.0022298, 0.0022233, 
    0.0022168, 0.0022105, 0.0022042, 0.0021979, 0.0021918, 0.0021856, 
    0.0021796, 0.0021736, 0.0021677, 0.0021619, 0.002156, 0.0021503, 
    0.0021445, 0.0021389, 0.0021332, 0.0021276, 0.0021221, 0.0021165, 
    0.002111, 0.0021056, 0.0021001, 0.0020947, 0.0020892, 0.0020838, 
    0.0020784, 0.002073, 0.0020676, 0.0020622, 0.0020568, 0.0020513, 
    0.0020459, 0.0020404, 0.0020349, 0.0020294, 0.0020238, 0.0020182, 
    0.0020126, 0.0020069, 0.0020012, 0.0019955, 0.0019897, 0.0019839, 
    0.001978, 0.0019721, 0.0019662, 0.0019602, 0.0019542, 0.0019481, 
    0.0019419, 0.0019358, 0.0019296, 0.0019233, 0.001917, 0.0019107, 
    0.0019043, 0.0018979, 0.0018915, 0.001885, 0.0018785, 0.001872, 
    0.0018655, 0.0018589, 0.0018523, 0.0018457, 0.001839, 0.0018324, 
    0.0018257, 0.0018191, 0.0018124, 0.0018057, 0.001799, 0.0017924, 
    0.0017857, 0.001779, 0.0017723, 0.0017656, 0.001759, 0.0017523, 
    0.0017456, 0.0017389, 0.0017323, 0.0017256, 0.0017189, 0.0017123, 
    0.0017057, 0.001699, 0.0016924, 0.0016859, 0.0016793, 0.0016728, 
    0.0016663, 0.0016599, 0.0016535, 0.0016472, 0.001641, 0.0016348, 
    0.0016286, 0.0016226, 0.0016166, 0.0016106, 0.0016048, 0.001599, 
    0.0015932, 0.0015875, 0.0015819, 0.0015763, 0.0015707, 0.0015651, 
    0.0015596, 0.001554, 0.0015485, 0.0015429, 0.0015374, 0.0015318, 
    0.0015262, 0.0015206, 0.001515, 0.0015097, 0.001504, 0.0014983, 
    0.0014926, 0.0014868, 0.0014811, 0.0014753, 0.0014696, 0.0014638, 
    0.001458, 0.0014523, 0.0014465, 0.0014408, 0.001435, 0.0014293, 
    0.0014236, 0.001418, 0.0014123, 0.0014066, 0.001401, 0.0013954, 
    0.0013898, 0.0013842, 0.0013786, 0.0013731, 0.0013675, 0.001362, 
    0.0013564, 0.0013509, 0.0013454, 0.0013399, 0.0013345, 0.001329, 
    0.0013236, 0.0013183, 0.001313, 0.0013077, 0.0013025, 0.0012974, 
    0.0012923, 0.0012873, 0.0012823, 0.0012774, 0.0012726, 0.0012678, 
    0.0012631, 0.0012585, 0.0012538, 0.0012493, 0.0012447, 0.0012402, 
    0.0012358, 0.0012313, 0.0012268, 0.0012224, 0.001218, 0.0012135, 
    0.001209, 0.0012046, 0.0012001, 0.0011955, 0.0011909, 0.0011863, 
    0.0011817, 0.0011769, 0.0011722, 0.0011674, 0.0011625, 0.0011575, 
    0.0011525, 0.0011475, 0.0011424, 0.0011372, 0.001132, 0.0011267, 
    0.0011213, 0.0011159, 0.0011105, 0.0011051, 0.0010996, 0.0010941, 
    0.0010886, 0.0010831, 0.0010776, 0.0010722, 0.0010668, 0.0010614, 
    0.0010561, 0.0010509, 0.0010458, 0.0010407, 0.0010357, 0.0010308, 
    0.0010261, 0.0010214, 0.0010168, 0.0010124, 0.001008, 0.0010037, 
    0.00099956, 0.00099548, 0.00099149, 0.00098759, 0.00098375, 0.00097998, 
    0.00097627, 0.00097262, 0.000969, 0.00096542, 0.00096187, 0.00095833, 
    0.00095481, 0.00095129, 0.00094777, 0.00094425, 0.00094071, 0.00093717, 
    0.00093361, 0.00093004, 0.00092645, 0.00092284, 0.00091922, 0.0009156, 
    0.00091196, 0.00090832, 0.00090467, 0.00090102, 0.00089738, 0.00089373, 
    0.00089008, 0.00088643, 0.00088278, 0.00087912, 0.00087545, 0.00087177, 
    0.00086807, 0.00086435, 0.0008606, 0.00085682, 0.00085299, 0.00084912, 
    0.0008452, 0.00084123, 0.00083721, 0.00083313, 0.00082899, 0.00082479, 
    0.00082055, 0.00081625, 0.00081191, 0.00080753, 0.00080312, 0.00079868, 
    0.00079422, 0.00078975, 0.00078528, 0.00078081, 0.00077636, 0.00077192, 
    0.00076751, 0.00076314, 0.0007588, 0.0007545, 0.00075025, 0.00074605, 
    0.0007419, 0.00073781, 0.00073378, 0.00072981, 0.0007259, 0.00072205, 
    0.00071827, 0.00071456, 0.00071092, 0.00070734, 0.00070384, 0.00070041, 
    0.00069705, 0.00069376, 0.00069054, 0.00068739, 0.0006843, 0.00068128, 
    0.00067831, 0.00067539, 0.00067253, 0.0006697, 0.00066691, 0.00066414, 
    0.0006614, 0.00065867, 0.00065595, 0.00065324, 0.00065053, 0.00064782, 
    0.0006451, 0.00064237, 0.00063964, 0.0006369, 0.00063414, 0.00063138, 
    0.00062861, 0.00062584, 0.00062305, 0.00062025, 0.00061745, 0.00061464, 
    0.00061182, 0.00060898, 0.00060614, 0.00060328, 0.0006004, 0.00059751, 
    0.00059461, 0.00059169, 0.00058875, 0.00058579, 0.00058283, 0.00057985, 
    0.00057686, 0.00057386, 0.00057087, 0.00056786, 0.00056486, 0.00056187, 
    0.00055888, 0.00055589, 0.00055291, 0.00054992, 0.00054694, 0.00054396, 
    0.00054098, 0.00053798, 0.00053497, 0.00053194, 0.00052889, 0.00052581, 
    0.0005227, 0.00051955, 0.00051638, 0.00051317, 0.00050994, 0.00050668, 
    0.00050339, 0.00050009, 0.00049679, 0.00049348, 0.00049018, 0.00048689, 
    0.00048363, 0.00048039, 0.0004772, 0.00047405, 0.00047096, 0.00046792, 
    0.00046495, 0.00046204, 0.0004592, 0.00045643, 0.00045375, 0.00045114, 
    0.00044861, 0.00044616, 0.00044379, 0.00044151, 0.0004393, 0.00043718, 
    0.00043514, 0.00043317, 0.00043127, 0.00042945, 0.00042769, 0.00042599, 
    0.00042435, 0.00042276, 0.0004212, 0.00041968, 0.00041819, 0.00041671, 
    0.00041525, 0.00041378, 0.00041231, 0.00041083, 0.00040933, 0.0004078, 
    0.00040624, 0.00040465, 0.00040302, 0.00040136, 0.00039965, 0.0003979, 
    0.00039611, 0.00039428, 0.00039241, 0.00039051, 0.00038857, 0.0003866, 
    0.0003846, 0.00038257, 0.00038052, 0.00037845, 0.00037635, 0.00037424, 
    0.00037212, 0.00036998, 0.00036784, 0.00036568, 0.00036353, 0.00036136, 
    0.0003592, 0.00035704, 0.00035488, 0.00035272, 0.00035057, 0.00034843, 
    0.00034629, 0.00034416, 0.00034205, 0.00033994, 0.00033784, 0.00033575, 
    0.00033368, 0.00033161, 0.00032955, 0.0003275, 0.00032546, 0.00032343, 
    0.0003214, 0.00031938, 0.00031737, 0.00031535, 0.00031335, 0.00031134, 
    0.00030934, 0.00030733, 0.00030533, 0.00030332, 0.00030131, 0.0002993, 
    0.00029728, 0.00029526, 0.00029323, 0.00029119, 0.00028914, 0.00028709, 
    0.00028503, 0.00028296, 0.00028089, 0.00027883, 0.00027676, 0.00027469, 
    0.00027264, 0.0002706, 0.00026857, 0.00026657, 0.00026459, 0.00026265, 
    0.00026073, 0.00025886, 0.00025703, 0.00025524, 0.0002535, 0.0002518, 
    0.00025016, 0.00024856, 0.00024702, 0.00024552, 0.00024407, 0.00024267, 
    0.0002413, 0.00023997, 0.00023868, 0.00023741, 0.00023617, 0.00023495, 
    0.00023374, 0.00023254, 0.00023135, 0.00023017, 0.00022898, 0.00022779, 
    0.0002266, 0.0002254, 0.00022418, 0.00022296, 0.00022172, 0.00022048, 
    0.00021921, 0.00021794, 0.00021666, 0.00021536, 0.00021405, 0.00021273, 
    0.0002114, 0.00021006, 0.00020872, 0.00020737, 0.00020601, 0.00020466, 
    0.00020331, 0.00020196, 0.00020062, 0.00019929, 0.00019797, 0.00019666, 
    0.00019536, 0.00019409, 0.00019283, 0.0001916, 0.00019039, 0.00018921, 
    0.00018804, 0.00018691, 0.00018579, 0.0001847, 0.00018363, 0.00018258, 
    0.00018156, 0.00018054, 0.00017954, 0.00017855, 0.00017758, 0.0001766, 
    0.00017564, 0.00017468, 0.00017372, 0.00017276, 0.00017181, 0.00017085, 
    0.0001699, 0.00016895, 0.00016799, 0.00016705, 0.0001661, 0.00016516, 
    0.00016423, 0.0001633, 0.00016238, 0.00016147, 0.00016058, 0.00015969, 
    0.00015882, 0.00015796, 0.00015711, 0.00015628, 0.00015546, 0.00015466, 
    0.00015386, 0.00015308, 0.00015231, 0.00015154, 0.00015078, 0.00015003, 
    0.00014929, 0.00014854, 0.0001478, 0.00014706, 0.00014632, 0.00014557, 
    0.00014482, 0.00014406, 0.00014329, 0.00014252, 0.00014174, 0.00014094, 
    0.00014014, 0.00013932, 0.00013849, 0.00013766, 0.00013681, 0.00013595, 
    0.00013508, 0.00013421, 0.00013333, 0.00013244, 0.00013155, 0.00013065, 
    0.00012976, 0.00012886, 0.00012796, 0.00012706, 0.00012617, 0.00012527, 
    0.00012438, 0.00012349, 0.0001226, 0.00012172, 0.00012084, 0.00011997, 
    0.0001191, 0.00011824, 0.00011739, 0.00011654, 0.0001157, 0.00011487, 
    0.00011406, 0.00011325, 0.00011246, 0.00011168, 0.00011092, 0.00011017, 
    0.00010943, 0.00010872, 0.00010802, 0.00010733, 0.00010666, 0.00010601, 
    0.00010536, 0.00010473, 0.00010411, 0.0001035, 0.00010289, 0.00010228, 
    0.00010168, 0.00010107, 0.00010046, 9.9851e-05, 9.9235e-05, 9.8614e-05, 
    9.7987e-05, 9.7354e-05, 9.6719e-05, 9.608e-05, 9.5441e-05, 9.48e-05, 
    9.4164e-05, 9.353e-05, 9.2904e-05, 9.2285e-05, 9.1678e-05, 9.1081e-05, 
    9.0499e-05, 8.9929e-05, 8.9377e-05, 8.8837e-05, 8.8316e-05, 8.7808e-05, 
    8.7317e-05, 8.6839e-05, 8.6374e-05, 8.5922e-05, 8.548e-05, 8.5047e-05, 
    8.4623e-05, 8.4204e-05, 8.3792e-05, 8.338e-05, 8.2973e-05, 8.2565e-05, 
    8.2156e-05, 8.1745e-05, 8.133e-05, 8.0912e-05, 8.0488e-05, 8.0059e-05, 
    7.9622e-05, 7.9179e-05, 7.8727e-05, 7.8268e-05, 7.78e-05, 7.7324e-05, 
    7.684e-05, 7.6346e-05, 7.5846e-05, 7.5338e-05, 7.4824e-05, 7.4302e-05, 
    7.3775e-05, 7.3243e-05, 7.2706e-05, 7.2167e-05, 7.1626e-05, 7.1083e-05, 
    7.0541e-05, 7e-05, 6.9461e-05, 6.8926e-05, 6.8395e-05, 6.787e-05, 
    6.7352e-05, 6.6842e-05, 6.6339e-05, 6.5846e-05, 6.5363e-05, 6.4891e-05, 
    6.4428e-05, 6.3979e-05, 6.3541e-05, 6.3115e-05, 6.2701e-05, 6.2299e-05, 
    6.191e-05, 6.1532e-05, 6.1167e-05, 6.0813e-05, 6.047e-05, 6.0137e-05, 
    5.9814e-05, 5.9499e-05, 5.9193e-05, 5.8894e-05, 5.8602e-05, 5.8315e-05, 
    5.8031e-05, 5.7752e-05, 5.7474e-05, 5.7198e-05, 5.6923e-05, 5.6646e-05, 
    5.637e-05, 5.6091e-05, 5.5812e-05, 5.5529e-05, 5.5244e-05, 5.4956e-05, 
    5.4666e-05, 5.4372e-05, 5.4077e-05, 5.3778e-05, 5.3478e-05, 5.3175e-05, 
    5.2871e-05, 5.2566e-05, 5.2259e-05, 5.1952e-05, 5.1644e-05, 5.1335e-05, 
    5.1026e-05, 5.0717e-05, 5.0408e-05, 5.0099e-05, 4.9789e-05, 4.948e-05, 
    4.9171e-05, 4.8862e-05, 4.8553e-05, 4.8245e-05, 4.7937e-05, 4.7631e-05, 
    4.7325e-05, 4.702e-05, 4.6717e-05, 4.6414e-05, 4.6114e-05, 4.5816e-05, 
    4.552e-05, 4.5226e-05, 4.4934e-05, 4.4646e-05, 4.436e-05, 4.4077e-05, 
    4.3796e-05, 4.3519e-05, 4.3245e-05, 4.2973e-05, 4.2704e-05, 4.2437e-05, 
    4.2174e-05, 4.1912e-05, 4.1653e-05, 4.1396e-05, 4.114e-05, 4.0888e-05, 
    4.0636e-05, 4.0387e-05, 4.0139e-05, 3.9894e-05, 3.965e-05, 3.9408e-05, 
    3.9168e-05, 3.893e-05, 3.8694e-05, 3.846e-05, 3.8229e-05, 3.7999e-05, 
    3.7772e-05, 3.7547e-05, 3.7324e-05, 3.7103e-05, 3.6884e-05, 3.6666e-05, 
    3.6451e-05, 3.6237e-05, 3.6023e-05, 3.5812e-05, 3.5601e-05, 3.5391e-05, 
    3.5181e-05, 3.4973e-05, 3.4765e-05, 3.4558e-05, 3.4351e-05, 3.4145e-05, 
    3.3939e-05, 3.3734e-05, 3.353e-05, 3.3326e-05, 3.3123e-05, 3.2921e-05, 
    3.272e-05, 3.2518e-05, 3.2318e-05, 3.2119e-05, 3.192e-05, 3.1722e-05, 
    3.1524e-05, 3.1327e-05, 3.1131e-05, 3.0936e-05, 3.0741e-05, 3.0548e-05, 
    3.0355e-05, 3.0164e-05, 2.9974e-05, 2.9785e-05, 2.9598e-05, 2.9412e-05, 
    2.9228e-05, 2.9046e-05, 2.8865e-05, 2.8687e-05, 2.851e-05, 2.8336e-05, 
    2.8163e-05, 2.7993e-05, 2.7825e-05, 2.7659e-05, 2.7494e-05, 2.7332e-05, 
    2.7171e-05, 2.7013e-05, 2.6856e-05, 2.67e-05, 2.6546e-05, 2.6394e-05, 
    2.6243e-05, 2.6093e-05, 2.5944e-05, 2.5797e-05, 2.565e-05, 2.5505e-05, 
    2.536e-05, 2.5216e-05, 2.5074e-05, 2.4932e-05, 2.479e-05, 2.465e-05, 
    2.451e-05, 2.437e-05, 2.4232e-05, 2.4094e-05, 2.3956e-05, 2.3819e-05, 
    2.3682e-05, 2.3545e-05, 2.3409e-05, 2.3273e-05, 2.3138e-05, 2.3004e-05, 
    2.287e-05, 2.2737e-05, 2.2604e-05, 2.2473e-05, 2.2343e-05, 2.2214e-05, 
    2.2086e-05, 2.196e-05, 2.1835e-05, 2.1713e-05, 2.1592e-05, 2.1473e-05, 
    2.1356e-05, 2.1241e-05, 2.1127e-05, 2.1016e-05, 2.0906e-05, 2.0798e-05, 
    2.0691e-05, 2.0585e-05, 2.048e-05, 2.0376e-05, 2.0272e-05, 2.0168e-05, 
    2.0065e-05, 1.996e-05, 1.9856e-05, 1.975e-05, 1.9644e-05, 1.9537e-05, 
    1.9429e-05, 1.932e-05, 1.921e-05, 1.9099e-05, 1.8987e-05, 1.8874e-05, 
    1.8761e-05, 1.8648e-05, 1.8535e-05, 1.8421e-05, 1.8308e-05, 1.8195e-05, 
    1.8083e-05, 1.7971e-05, 1.786e-05, 1.775e-05, 1.7641e-05, 1.7534e-05, 
    1.7427e-05, 1.7322e-05, 1.7219e-05, 1.7117e-05, 1.7017e-05, 1.6918e-05, 
    1.6822e-05, 1.6727e-05, 1.6633e-05, 1.6542e-05, 1.6452e-05, 1.6364e-05, 
    1.6277e-05, 1.6192e-05, 1.6108e-05, 1.6025e-05, 1.5944e-05, 1.5863e-05, 
    1.5784e-05, 1.5705e-05, 1.5627e-05, 1.5549e-05, 1.5472e-05, 1.5395e-05, 
    1.5318e-05, 1.5241e-05, 1.5164e-05, 1.5087e-05, 1.501e-05, 1.4933e-05, 
    1.4856e-05, 1.4778e-05, 1.47e-05, 1.4622e-05, 1.4544e-05, 1.4465e-05, 
    1.4386e-05, 1.4307e-05, 1.4228e-05, 1.4148e-05, 1.4069e-05, 1.3989e-05, 
    1.391e-05, 1.3831e-05, 1.3751e-05, 1.3673e-05, 1.3594e-05, 1.3516e-05, 
    1.3438e-05, 1.3361e-05, 1.3285e-05, 1.3209e-05, 1.3133e-05, 1.3058e-05, 
    1.2984e-05, 1.291e-05, 1.2837e-05, 1.2765e-05, 1.2693e-05, 1.2622e-05, 
    1.2551e-05, 1.2481e-05, 1.2411e-05, 1.2342e-05, 1.2274e-05, 1.2206e-05, 
    1.2138e-05, 1.2071e-05, 1.2005e-05, 1.1939e-05, 1.1873e-05, 1.1809e-05, 
    1.1744e-05, 1.1681e-05, 1.1617e-05, 1.1555e-05, 1.1493e-05, 1.1432e-05, 
    1.1371e-05, 1.1311e-05, 1.1252e-05, 1.1208e-05, 1.1164e-05, 1.1121e-05, 
    1.1079e-05, 1.1037e-05, 1.0996e-05, 1.0955e-05, 1.0914e-05, 1.0874e-05, 
    1.0834e-05, 1.0794e-05, 1.0754e-05, 1.0715e-05, 1.0676e-05, 1.0637e-05, 
    1.0598e-05, 1.0559e-05, 1.052e-05, 1.0481e-05, 1.0442e-05, 1.0404e-05, 
    1.0365e-05, 1.0326e-05, 1.0288e-05, 1.0249e-05, 1.0211e-05, 1.0172e-05, 
    1.0134e-05, 1.0096e-05, 1.0058e-05, 1.002e-05, 9.9825e-06, 9.945e-06, 
    9.9076e-06, 9.8704e-06, 9.8333e-06, 9.7964e-06, 9.7597e-06, 9.7231e-06, 
    9.6866e-06, 9.6502e-06, 9.6139e-06, 9.5777e-06, 9.5417e-06, 9.5056e-06, 
    9.4697e-06, 9.4338e-06, 9.398e-06, 9.3622e-06, 9.3265e-06, 9.2909e-06, 
    9.2554e-06, 9.2199e-06, 9.1846e-06, 9.1494e-06, 9.1144e-06, 9.0795e-06, 
    9.0448e-06, 9.0103e-06, 8.976e-06, 8.9419e-06, 8.9081e-06, 8.8744e-06, 
    8.8409e-06, 8.8077e-06, 8.7747e-06, 8.7419e-06, 8.7093e-06, 8.6769e-06, 
    8.6446e-06, 8.6124e-06, 8.5804e-06, 8.5486e-06, 8.5168e-06, 8.4851e-06, 
    8.4535e-06, 8.422e-06, 8.3906e-06, 8.3593e-06, 8.3281e-06, 8.2969e-06, 
    8.2659e-06, 8.235e-06, 8.2042e-06, 8.1735e-06, 8.143e-06, 8.1127e-06, 
    8.0825e-06, 8.0525e-06, 8.0227e-06, 7.9931e-06, 7.9636e-06, 7.9344e-06, 
    7.9052e-06, 7.8763e-06, 7.8476e-06, 7.8189e-06, 7.7905e-06, 7.7622e-06, 
    7.734e-06, 7.7059e-06, 7.678e-06, 7.6502e-06, 7.6225e-06, 7.5949e-06, 
    7.5674e-06, 7.54e-06, 7.5128e-06, 7.4857e-06, 7.4587e-06, 7.4319e-06, 
    7.4052e-06, 7.3787e-06, 7.3523e-06, 7.3261e-06, 7.3e-06, 7.2741e-06, 
    7.2483e-06, 7.2227e-06, 7.1972e-06, 7.1718e-06, 7.1465e-06, 7.1213e-06, 
    7.0962e-06, 7.0712e-06, 7.0462e-06, 7.0213e-06, 6.9964e-06, 6.9716e-06, 
    6.9467e-06, 6.922e-06, 6.8972e-06, 6.8725e-06, 6.8479e-06, 6.8232e-06, 
    6.7987e-06, 6.7742e-06, 6.7497e-06, 6.7254e-06, 6.7011e-06, 6.6768e-06, 
    6.6527e-06, 6.6286e-06, 6.6047e-06, 6.5808e-06, 6.557e-06, 6.5333e-06, 
    6.5097e-06, 6.4862e-06, 6.4628e-06, 6.4395e-06, 6.4163e-06, 6.3932e-06, 
    6.3701e-06, 6.3472e-06, 6.3243e-06, 6.3016e-06, 6.2789e-06, 6.2563e-06, 
    6.2338e-06, 6.2113e-06, 6.189e-06, 6.1667e-06, 6.1446e-06, 6.1225e-06, 
    6.1005e-06, 6.0786e-06, 6.0568e-06, 6.0351e-06, 6.0135e-06, 5.992e-06, 
    5.9705e-06, 5.9492e-06, 5.9279e-06, 5.9067e-06, 5.8856e-06, 5.8646e-06, 
    5.8437e-06, 5.8229e-06, 5.8021e-06, 5.7814e-06, 5.7608e-06, 5.7403e-06, 
    5.7198e-06, 5.6995e-06, 5.6792e-06, 5.6589e-06, 5.6388e-06, 5.6187e-06, 
    5.5987e-06, 5.5787e-06, 5.5589e-06, 5.5391e-06, 5.5194e-06, 5.4998e-06, 
    5.4803e-06, 5.4608e-06, 5.4415e-06, 5.4222e-06, 5.4031e-06, 5.384e-06, 
    5.3651e-06, 5.3463e-06, 5.3276e-06, 5.309e-06, 5.2905e-06, 5.2721e-06, 
    5.2538e-06, 5.2356e-06, 5.2176e-06, 5.1996e-06, 5.1817e-06, 5.1639e-06, 
    5.1462e-06, 5.1285e-06, 5.1109e-06, 5.0934e-06, 5.0759e-06, 5.0585e-06, 
    5.0411e-06, 5.0237e-06, 5.0063e-06, 4.989e-06, 4.9717e-06, 4.9545e-06, 
    4.9372e-06, 4.92e-06, 4.9029e-06, 4.8857e-06, 4.8686e-06, 4.8516e-06, 
    4.8346e-06, 4.8176e-06, 4.8007e-06, 4.7839e-06, 4.7671e-06, 4.7503e-06, 
    4.7337e-06, 4.7171e-06, 4.7005e-06, 4.6841e-06, 4.6677e-06, 4.6513e-06, 
    4.6351e-06, 4.6189e-06, 4.6027e-06, 4.5867e-06, 4.5707e-06, 4.5547e-06, 
    4.5388e-06, 4.523e-06, 4.5072e-06, 4.4915e-06, 4.4759e-06, 4.4603e-06, 
    4.4448e-06, 4.4293e-06, 4.4139e-06, 4.3985e-06, 4.3832e-06, 4.368e-06, 
    4.3528e-06, 4.3377e-06, 4.3226e-06, 4.3076e-06, 4.2926e-06, 4.2777e-06, 
    4.2629e-06, 4.2481e-06, 4.2334e-06, 4.2187e-06, 4.2041e-06, 4.1896e-06, 
    4.1751e-06, 4.1607e-06, 4.1463e-06, 4.132e-06, 4.1178e-06, 4.1036e-06, 
    4.0895e-06, 4.0754e-06, 4.0614e-06, 4.0474e-06, 4.0335e-06, 4.0196e-06, 
    4.0058e-06, 3.992e-06, 3.9783e-06, 3.9646e-06, 3.951e-06, 3.9374e-06, 
    3.9238e-06 ;

 bangle_L1_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_L2_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_sigma =
  0.00134, 0.0013437, 0.0013472, 0.0013502, 0.0013528, 0.0013553, 0.0013573, 
    0.0013592, 0.0013606, 0.0013618, 0.0013628, 0.0013638, 0.0013647, 
    0.0013655, 0.0013662, 0.0013668, 0.0013673, 0.0013676, 0.0013676, 
    0.0013673, 0.0013668, 0.001366, 0.0013652, 0.0013643, 0.0013634, 
    0.0013624, 0.0013616, 0.0013608, 0.0013603, 0.0013599, 0.0013597, 
    0.0013598, 0.0013601, 0.0013607, 0.0013615, 0.0013625, 0.0013636, 
    0.0013649, 0.0013663, 0.0013677, 0.0013691, 0.0013704, 0.0013716, 
    0.0013726, 0.0013735, 0.0013743, 0.0013749, 0.0013755, 0.001376, 
    0.0013765, 0.001377, 0.0013775, 0.0013781, 0.0013786, 0.0013792, 
    0.0013798, 0.0013805, 0.0013811, 0.0013818, 0.0013824, 0.0013831, 
    0.0013838, 0.0013845, 0.001385, 0.0013855, 0.001386, 0.0013865, 
    0.0013871, 0.0013877, 0.0013883, 0.001389, 0.0013898, 0.0013906, 
    0.0013915, 0.0013924, 0.0013933, 0.0013942, 0.001395, 0.0013956, 
    0.001396, 0.001396, 0.0013959, 0.0013956, 0.0013953, 0.0013949, 
    0.0013946, 0.0013943, 0.0013939, 0.0013934, 0.0013928, 0.0013922, 
    0.0013916, 0.0013911, 0.0013906, 0.0013902, 0.0013896, 0.0013891, 
    0.0013884, 0.0013878, 0.0013871, 0.0013865, 0.001386, 0.0013857, 
    0.0013854, 0.0013852, 0.0013851, 0.001385, 0.0013851, 0.0013852, 
    0.0013853, 0.0013852, 0.0013852, 0.0013849, 0.0013846, 0.0013842, 
    0.0013837, 0.0013832, 0.0013827, 0.0013821, 0.0013816, 0.0013811, 
    0.0013807, 0.0013804, 0.0013801, 0.0013799, 0.0013797, 0.0013796, 
    0.0013795, 0.0013795, 0.0013795, 0.0013795, 0.0013795, 0.0013796, 
    0.0013796, 0.0013797, 0.0013798, 0.0013799, 0.00138, 0.0013802, 
    0.0013803, 0.0013804, 0.0013804, 0.0013803, 0.0013802, 0.0013798, 
    0.0013792, 0.0013784, 0.0013771, 0.0013757, 0.001374, 0.0013722, 
    0.0013705, 0.0013691, 0.0013679, 0.0013671, 0.0013666, 0.0013664, 
    0.0013664, 0.0013667, 0.0013671, 0.0013675, 0.0013677, 0.0013677, 
    0.0013675, 0.0013665, 0.0013653, 0.001363, 0.00136, 0.0013562, 0.0013509, 
    0.0013451, 0.0013377, 0.0013293, 0.0013198, 0.0013088, 0.0012971, 
    0.001284, 0.0012702, 0.0012555, 0.0012398, 0.0012235, 0.0012061, 
    0.0011881, 0.0011692, 0.0011493, 0.0011287, 0.0011067, 0.0010843, 
    0.0010614, 0.0010386, 0.0010157, 0.0009934, 0.00097129, 0.00095024, 
    0.00093045, 0.0009114, 0.00089528, 0.00088002, 0.00086727, 0.0008562, 
    0.00084648, 0.00083964, 0.00083371, 0.00082995, 0.00082722, 0.00082546, 
    0.00082474, 0.00082431, 0.00082429, 0.00082424, 0.00082417, 0.00082376, 
    0.00082321, 0.00082216, 0.00082093, 0.00081946, 0.00081761, 0.0008156, 
    0.00081304, 0.00081032, 0.00080734, 0.00080406, 0.00080064, 0.00079656, 
    0.00079224, 0.00078745, 0.0007822, 0.00077669, 0.0007708, 0.00076483, 
    0.00075876, 0.00075272, 0.0007467, 0.00074081, 0.00073502, 0.00072958, 
    0.00072453, 0.00071978, 0.00071565, 0.0007117, 0.00070818, 0.00070493, 
    0.00070195, 0.00069941, 0.00069702, 0.00069506, 0.00069329, 0.00069174, 
    0.00069044, 0.00068923, 0.00068813, 0.00068708, 0.00068611, 0.00068523, 
    0.00068439, 0.00068375, 0.00068319, 0.00068276, 0.00068241, 0.00068211, 
    0.00068191, 0.00068175, 0.00068167, 0.00068165, 0.00068165, 0.00068167, 
    0.00068169, 0.00068171, 0.00068173, 0.00068175, 0.00068176, 0.00068177, 
    0.00068176, 0.00068176, 0.00068177, 0.00068179, 0.0006818, 0.00068183, 
    0.00068185, 0.00068187, 0.0006819, 0.00068192, 0.00068193, 0.00068194, 
    0.00068194, 0.00068194, 0.00068192, 0.0006819, 0.00068186, 0.00068182, 
    0.00068175, 0.00068168, 0.00068161, 0.00068153, 0.00068144, 0.00068136, 
    0.00068128, 0.0006812, 0.00068112, 0.00068106, 0.00068101, 0.00068096, 
    0.00068093, 0.00068091, 0.00068089, 0.00068087, 0.00068087, 0.00068088, 
    0.00068089, 0.0006809, 0.00068091, 0.00068091, 0.00068091, 0.0006809, 
    0.00068088, 0.00068084, 0.0006808, 0.00068074, 0.00068067, 0.0006806, 
    0.00068052, 0.00068044, 0.00068036, 0.00068027, 0.00068018, 0.00068009, 
    0.00067999, 0.00067988, 0.00067978, 0.00067966, 0.00067953, 0.00067939, 
    0.00067923, 0.00067907, 0.0006789, 0.00067872, 0.00067852, 0.00067833, 
    0.00067814, 0.00067796, 0.00067778, 0.00067762, 0.00067746, 0.00067731, 
    0.0006772, 0.00067711, 0.00067706, 0.00067703, 0.00067701, 0.00067702, 
    0.00067704, 0.00067707, 0.00067709, 0.0006771, 0.00067708, 0.00067704, 
    0.00067695, 0.00067682, 0.00067664, 0.00067639, 0.00067609, 0.00067565, 
    0.00067511, 0.00067445, 0.00067361, 0.00067269, 0.00067149, 0.00067014, 
    0.00066856, 0.0006666, 0.00066446, 0.00066169, 0.00065865, 0.00065508, 
    0.00065079, 0.00064608, 0.00064012, 0.00063376, 0.0006266, 0.00061873, 
    0.00061035, 0.00060117, 0.00059183, 0.00058243, 0.00057345, 0.00056477, 
    0.00055684, 0.00054915, 0.00054229, 0.00053603, 0.00053035, 0.00052544, 
    0.0005207, 0.00051623, 0.00051195, 0.00050789, 0.00050418, 0.00050061, 
    0.00049752, 0.00049475, 0.00049243, 0.00049063, 0.00048905, 0.00048802, 
    0.00048721, 0.00048676, 0.00048659, 0.00048655, 0.00048655, 0.0004865, 
    0.00048638, 0.00048605, 0.00048561, 0.00048463, 0.00048339, 0.00048157, 
    0.00047919, 0.00047643, 0.00047281, 0.00046899, 0.00046482, 0.00046058, 
    0.00045627, 0.00045246, 0.00044884, 0.00044579, 0.00044307, 0.00044067, 
    0.00043878, 0.00043703, 0.00043552, 0.00043397, 0.00043236, 0.00043057, 
    0.00042874, 0.00042688, 0.00042494, 0.0004229, 0.00042078, 0.00041863, 
    0.00041639, 0.00041405, 0.00041153, 0.00040924, 0.00040704, 0.00040533, 
    0.0004036, 0.00040186, 0.00039992, 0.00039786, 0.00039561, 0.00039318, 
    0.00039034, 0.00038738, 0.00038433, 0.0003812, 0.00037799, 0.00037457, 
    0.00037099, 0.00036728, 0.00036334, 0.00035928, 0.00035497, 0.00035039, 
    0.00034554, 0.00034027, 0.00033478, 0.00032882, 0.00032271, 0.00031644, 
    0.0003103, 0.00030417, 0.00029831, 0.00029244, 0.00028657, 0.00028117, 
    0.00027592, 0.0002714, 0.00026715, 0.00026338, 0.00026018, 0.00025721, 
    0.00025467, 0.00025223, 0.00025001, 0.00024806, 0.00024624, 0.00024501, 
    0.00024389, 0.00024302, 0.00024245, 0.00024208, 0.00024184, 0.00024163, 
    0.00024152, 0.00024142, 0.00024135, 0.00024129, 0.00024123, 0.00024117, 
    0.0002411, 0.00024101, 0.0002409, 0.00024077, 0.0002406, 0.00024039, 
    0.00024016, 0.00023987, 0.00023957, 0.0002392, 0.00023883, 0.00023846, 
    0.00023811, 0.00023776, 0.00023739, 0.00023697, 0.0002365, 0.00023592, 
    0.00023528, 0.00023427, 0.00023309, 0.00023159, 0.0002297, 0.00022759, 
    0.00022486, 0.00022188, 0.00021835, 0.0002143, 0.00020987, 0.0002047, 
    0.00019921, 0.00019315, 0.00018684, 0.00018028, 0.000174, 0.00016771, 
    0.0001618, 0.00015609, 0.00015058, 0.00014558, 0.00014069, 0.00013645, 
    0.00013247, 0.00012882, 0.00012557, 0.00012243, 0.0001197, 0.00011704, 
    0.00011454, 0.00011208, 0.00010961, 0.00010711, 0.00010461, 0.00010217, 
    9.9813e-05, 9.7464e-05, 9.5672e-05, 9.4122e-05, 9.3106e-05, 9.2456e-05, 
    9.2005e-05, 9.1868e-05, 9.1786e-05, 9.1811e-05, 9.1838e-05, 9.1864e-05, 
    9.1774e-05, 9.1625e-05, 9.1318e-05, 9.0887e-05, 9.0356e-05, 8.976e-05, 
    8.9151e-05, 8.854e-05, 8.7933e-05, 8.7332e-05, 8.6748e-05, 8.6168e-05, 
    8.5609e-05, 8.5067e-05, 8.4546e-05, 8.4056e-05, 8.3578e-05, 8.3165e-05, 
    8.2796e-05, 8.2489e-05, 8.2334e-05, 8.2254e-05, 8.2502e-05, 8.2862e-05, 
    8.3406e-05, 8.4089e-05, 8.483e-05, 8.5637e-05, 8.6394e-05, 8.7058e-05, 
    8.7603e-05, 8.8083e-05, 8.839e-05, 8.8647e-05, 8.8793e-05, 8.8869e-05, 
    8.89e-05, 8.8833e-05, 8.8753e-05, 8.8657e-05, 8.857e-05, 8.8489e-05, 
    8.8384e-05, 8.8273e-05, 8.8146e-05, 8.8032e-05, 8.793e-05, 8.7849e-05, 
    8.7772e-05, 8.7699e-05, 8.7606e-05, 8.749e-05, 8.7289e-05, 8.7052e-05, 
    8.6715e-05, 8.6359e-05, 8.5979e-05, 8.5613e-05, 8.5255e-05, 8.4961e-05, 
    8.4718e-05, 8.4562e-05, 8.4534e-05, 8.4564e-05, 8.4755e-05, 8.4977e-05, 
    8.5259e-05, 8.5517e-05, 8.5762e-05, 8.5954e-05, 8.6133e-05, 8.6287e-05, 
    8.6417e-05, 8.653e-05, 8.6585e-05, 8.6622e-05, 8.6618e-05, 8.6572e-05, 
    8.6494e-05, 8.635e-05, 8.6198e-05, 8.6054e-05, 8.5909e-05, 8.5762e-05, 
    8.5583e-05, 8.5403e-05, 8.5253e-05, 8.5128e-05, 8.5032e-05, 8.4931e-05, 
    8.4825e-05, 8.4681e-05, 8.4524e-05, 8.4349e-05, 8.4124e-05, 8.3878e-05, 
    8.3596e-05, 8.3301e-05, 8.2984e-05, 8.2612e-05, 8.2214e-05, 8.1778e-05, 
    8.1345e-05, 8.0924e-05, 8.0576e-05, 8.0266e-05, 8.0095e-05, 7.9954e-05, 
    7.9875e-05, 7.9831e-05, 7.981e-05, 7.9809e-05, 7.9804e-05, 7.9783e-05, 
    7.9747e-05, 7.9698e-05, 7.9626e-05, 7.9545e-05, 7.9442e-05, 7.9339e-05, 
    7.9234e-05, 7.9118e-05, 7.8997e-05, 7.8872e-05, 7.8763e-05, 7.8672e-05, 
    7.86e-05, 7.8531e-05, 7.8442e-05, 7.8342e-05, 7.8227e-05, 7.8095e-05, 
    7.7954e-05, 7.7776e-05, 7.7583e-05, 7.7368e-05, 7.7104e-05, 7.6817e-05, 
    7.6465e-05, 7.6112e-05, 7.5758e-05, 7.5415e-05, 7.5079e-05, 7.4796e-05, 
    7.4529e-05, 7.4299e-05, 7.4098e-05, 7.3918e-05, 7.3795e-05, 7.369e-05, 
    7.363e-05, 7.3584e-05, 7.3551e-05, 7.3516e-05, 7.3479e-05, 7.3435e-05, 
    7.3386e-05, 7.3331e-05, 7.3254e-05, 7.3161e-05, 7.3013e-05, 7.284e-05, 
    7.2639e-05, 7.2415e-05, 7.2182e-05, 7.1927e-05, 7.1664e-05, 7.139e-05, 
    7.1119e-05, 7.085e-05, 7.0607e-05, 7.0388e-05, 7.0209e-05, 7.0071e-05, 
    6.9951e-05, 6.9874e-05, 6.9806e-05, 6.9753e-05, 6.9718e-05, 6.9692e-05, 
    6.9681e-05, 6.9672e-05, 6.9669e-05, 6.9666e-05, 6.9666e-05, 6.9663e-05, 
    6.9657e-05, 6.9644e-05, 6.9627e-05, 6.9607e-05, 6.9587e-05, 6.9568e-05, 
    6.9547e-05, 6.9525e-05, 6.9501e-05, 6.9477e-05, 6.9456e-05, 6.9446e-05, 
    6.9442e-05, 6.9445e-05, 6.9448e-05, 6.9452e-05, 6.9456e-05, 6.9461e-05, 
    6.9466e-05, 6.9471e-05, 6.9476e-05, 6.9484e-05, 6.9492e-05, 6.9504e-05, 
    6.9509e-05, 6.9511e-05, 6.9504e-05, 6.9498e-05, 6.9497e-05, 6.95e-05, 
    6.9507e-05, 6.9511e-05, 6.9513e-05, 6.9513e-05, 6.9512e-05, 6.9511e-05, 
    6.951e-05, 6.9515e-05, 6.9537e-05, 6.9572e-05, 6.9617e-05, 6.9663e-05, 
    6.9709e-05, 6.9753e-05, 6.9799e-05, 6.9848e-05, 6.9896e-05, 6.9941e-05, 
    6.9971e-05, 7.0001e-05, 7.0028e-05, 7.0051e-05, 7.0074e-05, 7.0111e-05, 
    7.0153e-05, 7.02e-05, 7.0258e-05, 7.032e-05, 7.0391e-05, 7.046e-05, 
    7.0525e-05, 7.0579e-05, 7.0627e-05, 7.0659e-05, 7.0683e-05, 7.0694e-05, 
    7.069e-05, 7.0679e-05, 7.0656e-05, 7.0623e-05, 7.0567e-05, 7.0493e-05, 
    7.0407e-05, 7.0313e-05, 7.0218e-05, 7.0127e-05, 7.0038e-05, 6.995e-05, 
    6.9848e-05, 6.9735e-05, 6.9594e-05, 6.9428e-05, 6.9238e-05, 6.8996e-05, 
    6.8731e-05, 6.8397e-05, 6.8019e-05, 6.7591e-05, 6.7099e-05, 6.6586e-05, 
    6.6053e-05, 6.5539e-05, 6.5051e-05, 6.4599e-05, 6.4163e-05, 6.38e-05, 
    6.3466e-05, 6.318e-05, 6.2935e-05, 6.2709e-05, 6.2538e-05, 6.2381e-05, 
    6.2251e-05, 6.2132e-05, 6.2019e-05, 6.192e-05, 6.183e-05, 6.176e-05, 
    6.1708e-05, 6.1667e-05, 6.1644e-05, 6.1623e-05, 6.1609e-05, 6.1594e-05, 
    6.1578e-05, 6.1563e-05, 6.1549e-05, 6.1542e-05, 6.1539e-05, 6.154e-05, 
    6.154e-05, 6.1539e-05, 6.153e-05, 6.1511e-05, 6.148e-05, 6.1428e-05, 
    6.1367e-05, 6.1284e-05, 6.1197e-05, 6.1103e-05, 6.1003e-05, 6.0903e-05, 
    6.0816e-05, 6.0735e-05, 6.0662e-05, 6.0595e-05, 6.0531e-05, 6.0472e-05, 
    6.0415e-05, 6.036e-05, 6.0302e-05, 6.0242e-05, 6.0166e-05, 6.0089e-05, 
    6.0009e-05, 5.9926e-05, 5.9842e-05, 5.9752e-05, 5.9661e-05, 5.9567e-05, 
    5.9473e-05, 5.9378e-05, 5.9289e-05, 5.9205e-05, 5.914e-05, 5.9086e-05, 
    5.9044e-05, 5.9014e-05, 5.8989e-05, 5.8975e-05, 5.8964e-05, 5.8957e-05, 
    5.8954e-05, 5.8951e-05, 5.8951e-05, 5.8948e-05, 5.8944e-05, 5.8938e-05, 
    5.8932e-05, 5.8919e-05, 5.8902e-05, 5.8877e-05, 5.8841e-05, 5.8799e-05, 
    5.8737e-05, 5.8667e-05, 5.8583e-05, 5.8487e-05, 5.8386e-05, 5.827e-05, 
    5.8156e-05, 5.8047e-05, 5.7958e-05, 5.7881e-05, 5.7846e-05, 5.7822e-05, 
    5.7818e-05, 5.7815e-05, 5.7813e-05, 5.7792e-05, 5.7765e-05, 5.772e-05, 
    5.7669e-05, 5.7613e-05, 5.7553e-05, 5.7494e-05, 5.7447e-05, 5.7416e-05, 
    5.7401e-05, 5.7405e-05, 5.7415e-05, 5.7436e-05, 5.7458e-05, 5.748e-05, 
    5.7493e-05, 5.7503e-05, 5.7504e-05, 5.7506e-05, 5.7511e-05, 5.7522e-05, 
    5.7535e-05, 5.7516e-05, 5.7462e-05, 5.734e-05, 5.7114e-05, 5.6831e-05, 
    5.6318e-05, 5.5703e-05, 5.4859e-05, 5.3839e-05, 5.2692e-05, 5.1357e-05, 
    4.9968e-05, 4.8521e-05, 4.7193e-05, 4.5957e-05, 4.4988e-05, 4.4096e-05, 
    4.3422e-05, 4.2866e-05, 4.2426e-05, 4.2136e-05, 4.1894e-05, 4.1762e-05, 
    4.166e-05, 4.159e-05, 4.1539e-05, 4.1492e-05, 4.1439e-05, 4.1379e-05, 
    4.1306e-05, 4.118e-05, 4.1029e-05, 4.0787e-05, 4.0505e-05, 4.0158e-05, 
    3.9831e-05, 3.9515e-05, 3.9383e-05, 3.9307e-05, 3.9344e-05, 3.9457e-05, 
    3.9611e-05, 3.9786e-05, 3.9939e-05, 4.0037e-05, 4.0038e-05, 3.9978e-05, 
    3.972e-05, 3.9391e-05, 3.8885e-05, 3.8295e-05, 3.7634e-05, 3.701e-05, 
    3.6399e-05, 3.5855e-05, 3.5345e-05, 3.4869e-05, 3.4452e-05, 3.4058e-05, 
    3.3741e-05, 3.3469e-05, 3.3247e-05, 3.3074e-05, 3.292e-05, 3.2821e-05, 
    3.2746e-05, 3.2703e-05, 3.2682e-05, 3.2669e-05, 3.2665e-05, 3.2661e-05, 
    3.2659e-05, 3.2654e-05, 3.2647e-05, 3.2642e-05, 3.2642e-05, 3.2649e-05, 
    3.2662e-05, 3.2678e-05, 3.2695e-05, 3.2711e-05, 3.2724e-05, 3.274e-05, 
    3.2756e-05, 3.2778e-05, 3.28e-05, 3.282e-05, 3.2842e-05, 3.2866e-05, 
    3.2886e-05, 3.2905e-05, 3.2922e-05, 3.2937e-05, 3.295e-05, 3.2961e-05, 
    3.297e-05, 3.2973e-05, 3.2975e-05, 3.2976e-05, 3.2977e-05, 3.2977e-05, 
    3.2975e-05, 3.2973e-05, 3.2971e-05, 3.297e-05, 3.297e-05, 3.2972e-05, 
    3.2973e-05, 3.2975e-05, 3.2975e-05, 3.2974e-05, 3.2976e-05, 3.2977e-05, 
    3.2976e-05, 3.2962e-05, 3.2942e-05, 3.2908e-05, 3.2874e-05, 3.284e-05, 
    3.2818e-05, 3.2803e-05, 3.2805e-05, 3.2809e-05, 3.2819e-05, 3.283e-05, 
    3.2842e-05, 3.2866e-05, 3.2891e-05, 3.2919e-05, 3.2944e-05, 3.2965e-05, 
    3.2984e-05, 3.3005e-05, 3.3035e-05, 3.3059e-05, 3.3079e-05, 3.3093e-05, 
    3.3104e-05, 3.3115e-05, 3.3124e-05, 3.313e-05, 3.3135e-05, 3.3138e-05, 
    3.3146e-05, 3.3156e-05, 3.3169e-05, 3.3184e-05, 3.3202e-05, 3.3226e-05, 
    3.3251e-05, 3.3279e-05, 3.3306e-05, 3.3331e-05, 3.3356e-05, 3.3381e-05, 
    3.3407e-05, 3.3433e-05, 3.3458e-05, 3.3486e-05, 3.3513e-05, 3.3535e-05, 
    3.3553e-05, 3.3565e-05, 3.3564e-05, 3.356e-05, 3.3551e-05, 3.3544e-05, 
    3.3539e-05, 3.3537e-05, 3.3535e-05, 3.3529e-05, 3.3521e-05, 3.3512e-05, 
    3.3502e-05, 3.3492e-05, 3.3487e-05, 3.3484e-05, 3.3481e-05, 3.3483e-05, 
    3.3487e-05, 3.3496e-05, 3.3505e-05, 3.3514e-05, 3.3523e-05, 3.3533e-05, 
    3.3548e-05, 3.3566e-05, 3.359e-05, 3.3617e-05, 3.3647e-05, 3.369e-05, 
    3.3732e-05, 3.3767e-05, 3.3785e-05, 3.3792e-05, 3.38e-05, 3.381e-05, 
    3.3823e-05, 3.3823e-05, 3.3814e-05, 3.3786e-05, 3.3752e-05, 3.3707e-05, 
    3.3648e-05, 3.3578e-05, 3.3486e-05, 3.3389e-05, 3.3286e-05, 3.3171e-05, 
    3.3043e-05, 3.2895e-05, 3.2738e-05, 3.2562e-05, 3.2377e-05, 3.2183e-05, 
    3.1978e-05, 3.177e-05, 3.1566e-05, 3.1377e-05, 3.1213e-05, 3.1052e-05, 
    3.0892e-05, 3.0741e-05, 3.0588e-05, 3.0433e-05, 3.029e-05, 3.0154e-05, 
    3.0007e-05, 2.9854e-05, 2.9686e-05, 2.9524e-05, 2.9366e-05, 2.9234e-05, 
    2.9105e-05, 2.8982e-05, 2.8874e-05, 2.8778e-05, 2.8726e-05, 2.8685e-05, 
    2.8666e-05, 2.8662e-05, 2.8673e-05, 2.871e-05, 2.8757e-05, 2.8819e-05, 
    2.8878e-05, 2.8931e-05, 2.8984e-05, 2.9037e-05, 2.9083e-05, 2.9114e-05, 
    2.9125e-05, 2.9102e-05, 2.9065e-05, 2.9007e-05, 2.8944e-05, 2.887e-05, 
    2.8792e-05, 2.871e-05, 2.8619e-05, 2.8529e-05, 2.844e-05, 2.8364e-05, 
    2.8296e-05, 2.8244e-05, 2.8194e-05, 2.8149e-05, 2.8115e-05, 2.8088e-05, 
    2.8076e-05, 2.8067e-05, 2.8061e-05, 2.8061e-05, 2.8066e-05, 2.8074e-05, 
    2.8083e-05, 2.8097e-05, 2.811e-05, 2.8124e-05, 2.8144e-05, 2.8165e-05, 
    2.8185e-05, 2.8203e-05, 2.8218e-05, 2.8234e-05, 2.8251e-05, 2.8273e-05, 
    2.8294e-05, 2.8316e-05, 2.8342e-05, 2.837e-05, 2.8401e-05, 2.843e-05, 
    2.8456e-05, 2.8479e-05, 2.8499e-05, 2.8495e-05, 2.8487e-05, 2.8473e-05, 
    2.8451e-05, 2.8425e-05, 2.8404e-05, 2.8378e-05, 2.834e-05, 2.8308e-05, 
    2.8279e-05, 2.8257e-05, 2.8237e-05, 2.822e-05, 2.8203e-05, 2.8186e-05, 
    2.8168e-05, 2.815e-05, 2.8131e-05, 2.8115e-05, 2.8103e-05, 2.8097e-05, 
    2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8093e-05, 
    2.81e-05, 2.8111e-05, 2.8128e-05, 2.8147e-05, 2.8168e-05, 2.8215e-05, 
    2.8271e-05, 2.834e-05, 2.8425e-05, 2.8516e-05, 2.8617e-05, 2.8712e-05, 
    2.88e-05, 2.887e-05, 2.8931e-05, 2.8979e-05, 2.9025e-05, 2.9069e-05, 
    2.9106e-05, 2.9137e-05, 2.9163e-05, 2.9186e-05, 2.9206e-05, 2.9226e-05, 
    2.9245e-05, 2.9265e-05, 2.9286e-05, 2.9308e-05, 2.9328e-05, 2.9348e-05, 
    2.9366e-05, 2.9382e-05, 2.9396e-05, 2.9412e-05, 2.9431e-05, 2.9455e-05, 
    2.948e-05, 2.9504e-05, 2.9527e-05, 2.9548e-05, 2.9566e-05, 2.9583e-05, 
    2.9603e-05, 2.9622e-05, 2.9637e-05, 2.9653e-05, 2.967e-05, 2.9678e-05, 
    2.9683e-05, 2.9685e-05, 2.9688e-05, 2.969e-05, 2.9706e-05, 2.9722e-05, 
    2.9736e-05, 2.9753e-05, 2.9771e-05, 2.9795e-05, 2.982e-05, 2.9848e-05, 
    2.9878e-05, 2.991e-05, 2.9947e-05, 2.9987e-05, 3.0027e-05, 3.0064e-05, 
    3.0099e-05, 3.0126e-05, 3.0152e-05, 3.0173e-05, 3.0193e-05, 3.0212e-05, 
    3.0223e-05, 3.023e-05, 3.0226e-05, 3.0214e-05, 3.0193e-05, 3.0153e-05, 
    3.0105e-05, 3.0043e-05, 2.997e-05, 2.9881e-05, 2.9778e-05, 2.9669e-05, 
    2.954e-05, 2.9406e-05, 2.9264e-05, 2.9103e-05, 2.8933e-05, 2.8747e-05, 
    2.8548e-05, 2.8321e-05, 2.8073e-05, 2.781e-05, 2.7528e-05, 2.7246e-05, 
    2.6973e-05, 2.6698e-05, 2.6424e-05, 2.6148e-05, 2.5875e-05, 2.5614e-05, 
    2.5371e-05, 2.5144e-05, 2.4953e-05, 2.4774e-05, 2.4626e-05, 2.4484e-05, 
    2.435e-05, 2.4189e-05, 2.4022e-05, 2.3855e-05, 2.3698e-05, 2.3555e-05, 
    2.3427e-05, 2.3305e-05, 2.3202e-05, 2.3101e-05, 2.3001e-05, 2.2912e-05, 
    2.2828e-05, 2.2745e-05, 2.2667e-05, 2.2602e-05, 2.255e-05, 2.2505e-05, 
    2.2452e-05, 2.2401e-05, 2.2351e-05, 2.2313e-05, 2.2282e-05, 2.2258e-05, 
    2.2234e-05, 2.2208e-05, 2.2186e-05, 2.2166e-05, 2.2147e-05, 2.213e-05, 
    2.212e-05, 2.2115e-05, 2.2115e-05, 2.2113e-05, 2.211e-05, 2.2105e-05, 
    2.2104e-05, 2.2107e-05, 2.211e-05, 2.2113e-05, 2.2112e-05, 2.2111e-05, 
    2.2108e-05, 2.2108e-05, 2.2109e-05, 2.2109e-05, 2.2112e-05, 2.2117e-05, 
    2.2122e-05, 2.2125e-05, 2.2125e-05, 2.2125e-05, 2.2126e-05, 2.2125e-05, 
    2.2125e-05, 2.2125e-05, 2.2126e-05, 2.213e-05, 2.2139e-05, 2.2152e-05, 
    2.2176e-05, 2.2199e-05, 2.2217e-05, 2.2228e-05, 2.2234e-05, 2.2243e-05, 
    2.2253e-05, 2.2268e-05, 2.2283e-05, 2.2299e-05, 2.2313e-05, 2.2327e-05, 
    2.2339e-05, 2.2352e-05, 2.2366e-05, 2.2376e-05, 2.2382e-05, 2.2372e-05, 
    2.2355e-05, 2.2329e-05, 2.2298e-05, 2.2265e-05, 2.2227e-05, 2.2184e-05, 
    2.2134e-05, 2.2094e-05, 2.2059e-05, 2.2031e-05, 2.2002e-05, 2.1972e-05, 
    2.1947e-05, 2.1926e-05, 2.1913e-05, 2.1901e-05, 2.1887e-05, 2.187e-05, 
    2.185e-05, 2.1823e-05, 2.1795e-05, 2.1761e-05, 2.1728e-05, 2.1694e-05, 
    2.1667e-05, 2.1641e-05, 2.1616e-05, 2.1586e-05, 2.155e-05, 2.1509e-05, 
    2.1466e-05, 2.1427e-05, 2.1389e-05, 2.1355e-05, 2.1324e-05, 2.1295e-05, 
    2.1274e-05, 2.1257e-05, 2.1246e-05, 2.124e-05, 2.1236e-05, 2.1238e-05, 
    2.1243e-05, 2.1251e-05, 2.1262e-05, 2.1274e-05, 2.129e-05, 2.1305e-05, 
    2.1321e-05, 2.1339e-05, 2.1358e-05, 2.1377e-05, 2.1392e-05, 2.1397e-05, 
    2.1399e-05, 2.1398e-05, 2.1393e-05, 2.1385e-05, 2.1367e-05, 2.1343e-05, 
    2.1313e-05, 2.1272e-05, 2.1226e-05, 2.1162e-05, 2.1098e-05, 2.1031e-05, 
    2.098e-05, 2.0931e-05, 2.0875e-05, 2.0814e-05, 2.0747e-05, 2.0687e-05, 
    2.063e-05, 2.0594e-05, 2.0562e-05, 2.0535e-05, 2.0519e-05, 2.0507e-05, 
    2.0508e-05, 2.0505e-05, 2.0498e-05, 2.0484e-05, 2.0466e-05, 2.0439e-05, 
    2.0413e-05, 2.0386e-05, 2.035e-05, 2.0308e-05, 2.0288e-05, 2.0272e-05, 
    2.0263e-05, 2.0254e-05, 2.0245e-05, 2.0236e-05, 2.0228e-05, 2.0226e-05, 
    2.0235e-05, 2.0251e-05, 2.0297e-05, 2.0352e-05, 2.0429e-05, 2.0531e-05, 
    2.0656e-05, 2.0826e-05, 2.1016e-05, 2.1268e-05, 2.1561e-05, 2.1897e-05, 
    2.2239e-05, 2.2577e-05, 2.2895e-05, 2.3225e-05, 2.3571e-05, 2.3945e-05, 
    2.4323e-05, 2.4676e-05, 2.5003e-05, 2.5292e-05, 2.5555e-05, 2.5803e-05, 
    2.6005e-05, 2.6193e-05, 2.6352e-05, 2.6499e-05, 2.664e-05, 2.677e-05, 
    2.6892e-05, 2.6995e-05, 2.7091e-05, 2.7182e-05, 2.727e-05, 2.7354e-05, 
    2.7428e-05, 2.7495e-05, 2.7557e-05, 2.7599e-05, 2.7634e-05, 2.7653e-05, 
    2.7671e-05, 2.7688e-05, 2.7698e-05, 2.7707e-05, 2.7711e-05, 2.7718e-05, 
    2.7728e-05, 2.7738e-05, 2.7749e-05, 2.7765e-05, 2.7783e-05, 2.7802e-05, 
    2.7824e-05, 2.7846e-05, 2.786e-05, 2.7874e-05, 2.7887e-05, 2.7897e-05, 
    2.7905e-05, 2.7907e-05, 2.7905e-05, 2.7894e-05, 2.7882e-05, 2.7869e-05, 
    2.7847e-05, 2.782e-05, 2.7785e-05, 2.7749e-05, 2.7714e-05, 2.7682e-05, 
    2.7655e-05, 2.764e-05, 2.7631e-05, 2.7627e-05, 2.7628e-05, 2.763e-05, 
    2.7639e-05, 2.7654e-05, 2.7676e-05, 2.7712e-05, 2.7756e-05, 2.7818e-05, 
    2.789e-05, 2.7972e-05, 2.8074e-05, 2.8183e-05, 2.8306e-05, 2.8425e-05, 
    2.854e-05, 2.8642e-05, 2.8738e-05, 2.881e-05, 2.8874e-05, 2.8924e-05, 
    2.8962e-05, 2.8994e-05, 2.9014e-05, 2.9028e-05, 2.903e-05, 2.9021e-05, 
    2.9005e-05, 2.8987e-05, 2.8961e-05, 2.8918e-05, 2.8865e-05, 2.8805e-05, 
    2.8735e-05, 2.8666e-05, 2.8606e-05, 2.8567e-05, 2.8544e-05, 2.8571e-05, 
    2.8614e-05, 2.8693e-05, 2.879e-05, 2.8904e-05, 2.9042e-05, 2.9187e-05, 
    2.9344e-05, 2.9498e-05, 2.9651e-05, 2.9789e-05, 2.9922e-05, 3.0038e-05, 
    3.0143e-05, 3.0235e-05, 3.031e-05, 3.0378e-05, 3.0427e-05, 3.0469e-05, 
    3.0498e-05, 3.0512e-05, 3.0519e-05, 3.0509e-05, 3.0497e-05, 3.0479e-05, 
    3.0455e-05, 3.0428e-05, 3.0396e-05, 3.0361e-05, 3.0316e-05, 3.0274e-05, 
    3.0233e-05, 3.0186e-05, 3.0143e-05, 3.0109e-05, 3.0081e-05, 3.0056e-05, 
    3.0046e-05, 3.0039e-05, 3.0039e-05, 3.004e-05, 3.0043e-05, 3.0045e-05, 
    3.0046e-05, 3.0043e-05, 3.0037e-05, 3.0025e-05, 3.0004e-05, 2.9979e-05, 
    2.9948e-05, 2.9916e-05, 2.988e-05, 2.9847e-05, 2.9814e-05, 2.9788e-05, 
    2.9763e-05, 2.9738e-05, 2.9716e-05, 2.9695e-05, 2.9685e-05, 2.9677e-05, 
    2.9676e-05, 2.968e-05, 2.9688e-05, 2.9706e-05, 2.9726e-05, 2.9751e-05, 
    2.9782e-05, 2.9817e-05, 2.9856e-05, 2.9894e-05, 2.9928e-05, 2.9957e-05, 
    2.9982e-05, 2.9998e-05, 3.0013e-05, 3.0028e-05, 3.004e-05, 3.0048e-05, 
    3.0054e-05, 3.0058e-05, 3.0061e-05, 3.0062e-05, 3.0062e-05, 3.006e-05, 
    3.0057e-05, 3.0052e-05, 3.0045e-05, 3.0036e-05, 3.0022e-05, 3.0007e-05, 
    2.9987e-05, 2.9965e-05, 2.9938e-05, 2.9909e-05, 2.9879e-05, 2.9856e-05, 
    2.9837e-05, 2.9824e-05, 2.9814e-05, 2.9804e-05, 2.9796e-05, 2.9789e-05, 
    2.978e-05, 2.9779e-05, 2.9782e-05, 2.9801e-05, 2.9823e-05, 2.9854e-05, 
    2.9881e-05, 2.9905e-05, 2.9912e-05, 2.9916e-05, 2.992e-05, 2.9923e-05, 
    2.9925e-05, 2.9924e-05, 2.9921e-05, 2.9918e-05, 2.9918e-05, 2.9922e-05, 
    2.9928e-05, 2.9934e-05, 2.9938e-05, 2.9938e-05, 2.9935e-05, 2.993e-05, 
    2.9924e-05, 2.9916e-05, 2.9909e-05, 2.9904e-05, 2.9899e-05, 2.9894e-05, 
    2.9881e-05, 2.9872e-05, 2.9869e-05, 2.9872e-05, 2.9878e-05, 2.9892e-05, 
    2.9904e-05, 2.9913e-05, 2.9918e-05, 2.9921e-05, 2.9926e-05, 2.9932e-05, 
    2.9943e-05, 2.9958e-05, 2.9976e-05, 2.9986e-05, 2.9995e-05, 2.9997e-05, 
    2.9997e-05, 2.9993e-05, 2.9981e-05, 2.9968e-05, 2.9948e-05, 2.9932e-05, 
    2.992e-05, 2.9922e-05, 2.9929e-05, 2.9941e-05, 2.995e-05, 2.9956e-05, 
    2.9957e-05, 2.9957e-05, 2.996e-05, 2.9964e-05, 2.9969e-05, 2.9973e-05, 
    2.9977e-05, 2.9984e-05, 2.9989e-05, 2.9988e-05, 2.9991e-05, 2.9996e-05, 
    3.0011e-05, 3.0031e-05, 3.0063e-05, 3.0092e-05, 3.0121e-05, 3.0134e-05, 
    3.0144e-05, 3.0146e-05, 3.0146e-05, 3.0145e-05, 3.0143e-05, 3.0142e-05, 
    3.014e-05, 3.0141e-05, 3.0143e-05, 3.015e-05, 3.016e-05, 3.0175e-05, 
    3.0191e-05, 3.0208e-05, 3.0223e-05, 3.0236e-05, 3.0244e-05, 3.0251e-05, 
    3.0255e-05, 3.0257e-05, 3.0258e-05, 3.0256e-05, 3.0253e-05, 3.0249e-05, 
    3.0244e-05, 3.024e-05, 3.0244e-05, 3.0251e-05, 3.0267e-05, 3.0294e-05, 
    3.0325e-05, 3.0345e-05, 3.0365e-05, 3.0389e-05, 3.0419e-05, 3.0455e-05, 
    3.0504e-05, 3.0557e-05, 3.0615e-05, 3.0684e-05, 3.0761e-05, 3.0862e-05, 
    3.0971e-05, 3.1098e-05, 3.1242e-05, 3.14e-05, 3.1585e-05, 3.1777e-05, 
    3.1979e-05, 3.2181e-05, 3.2385e-05, 3.2562e-05, 3.2729e-05, 3.2876e-05, 
    3.3014e-05, 3.3138e-05, 3.3259e-05, 3.3378e-05, 3.3497e-05, 3.3616e-05, 
    3.3734e-05, 3.3837e-05, 3.3933e-05, 3.3999e-05, 3.4055e-05, 3.4092e-05, 
    3.4117e-05, 3.4136e-05, 3.4156e-05, 3.4179e-05, 3.4208e-05, 3.4225e-05, 
    3.4236e-05, 3.4237e-05, 3.4238e-05, 3.4239e-05, 3.4242e-05, 3.4247e-05, 
    3.4253e-05, 3.4258e-05, 3.4262e-05, 3.4265e-05, 3.4266e-05, 3.4265e-05, 
    3.4263e-05, 3.426e-05, 3.4255e-05, 3.4248e-05, 3.4235e-05, 3.4219e-05, 
    3.4188e-05, 3.4151e-05, 3.4106e-05, 3.404e-05, 3.3963e-05, 3.3853e-05, 
    3.3724e-05, 3.3562e-05, 3.3357e-05, 3.3132e-05, 3.2897e-05, 3.266e-05, 
    3.2425e-05, 3.2164e-05, 3.1889e-05, 3.1571e-05, 3.125e-05, 3.0926e-05, 
    3.0619e-05, 3.0322e-05, 3.0058e-05, 2.9802e-05, 2.9567e-05, 2.935e-05, 
    2.9146e-05, 2.8969e-05, 2.8801e-05, 2.8658e-05, 2.8529e-05, 2.8414e-05, 
    2.8318e-05, 2.8227e-05, 2.8142e-05, 2.8063e-05, 2.7989e-05, 2.7917e-05, 
    2.7847e-05, 2.7783e-05, 2.7725e-05, 2.7672e-05, 2.762e-05, 2.7569e-05, 
    2.7521e-05, 2.7471e-05, 2.7417e-05, 2.736e-05, 2.7302e-05, 2.7245e-05, 
    2.7189e-05, 2.7135e-05, 2.7078e-05, 2.7021e-05, 2.6967e-05, 2.6914e-05, 
    2.6866e-05, 2.6824e-05, 2.6785e-05, 2.6757e-05, 2.6732e-05, 2.6713e-05, 
    2.6697e-05, 2.6685e-05, 2.6675e-05, 2.6665e-05, 2.6658e-05, 2.6652e-05, 
    2.6647e-05, 2.6644e-05, 2.6641e-05, 2.664e-05, 2.6642e-05, 2.6649e-05, 
    2.6658e-05, 2.6669e-05, 2.6677e-05, 2.6684e-05, 2.6687e-05, 2.6686e-05, 
    2.6682e-05, 2.6656e-05, 2.6618e-05, 2.656e-05, 2.6479e-05, 2.6387e-05, 
    2.6269e-05, 2.6145e-05, 2.6011e-05, 2.5883e-05, 2.5759e-05, 2.5654e-05, 
    2.5559e-05, 2.5486e-05, 2.5433e-05, 2.5394e-05, 2.5385e-05, 2.5381e-05, 
    2.5387e-05, 2.5401e-05, 2.5421e-05, 2.5453e-05, 2.5488e-05, 2.553e-05, 
    2.5569e-05, 2.5606e-05, 2.5635e-05, 2.5661e-05, 2.5674e-05, 2.5681e-05, 
    2.5681e-05, 2.5658e-05, 2.5625e-05, 2.5558e-05, 2.5473e-05, 2.5366e-05, 
    2.5239e-05, 2.5105e-05, 2.4962e-05, 2.4813e-05, 2.4654e-05, 2.4487e-05, 
    2.4315e-05, 2.4147e-05, 2.3982e-05, 2.3827e-05, 2.3691e-05, 2.3566e-05, 
    2.348e-05, 2.3402e-05, 2.3342e-05, 2.3297e-05, 2.3262e-05, 2.324e-05, 
    2.3222e-05, 2.3211e-05, 2.3209e-05, 2.3212e-05, 2.3219e-05, 2.3227e-05, 
    2.3232e-05, 2.3236e-05, 2.3237e-05, 2.3236e-05, 2.3233e-05, 2.3227e-05, 
    2.3217e-05, 2.3202e-05, 2.3178e-05, 2.3148e-05, 2.31e-05, 2.3046e-05, 
    2.2981e-05, 2.2914e-05, 2.2845e-05, 2.2779e-05, 2.2717e-05, 2.2662e-05, 
    2.2623e-05, 2.259e-05, 2.2585e-05, 2.2587e-05, 2.2603e-05, 2.2624e-05, 
    2.2648e-05, 2.2664e-05, 2.2676e-05, 2.268e-05, 2.2682e-05, 2.2682e-05, 
    2.2682e-05, 2.2683e-05, 2.2688e-05, 2.2701e-05, 2.2719e-05, 2.2744e-05, 
    2.2767e-05, 2.2781e-05, 2.2782e-05, 2.2773e-05, 2.274e-05, 2.27e-05, 
    2.2648e-05, 2.26e-05, 2.2555e-05, 2.2517e-05, 2.2482e-05, 2.2461e-05, 
    2.2439e-05, 2.2416e-05, 2.2401e-05, 2.2389e-05, 2.2383e-05, 2.238e-05, 
    2.238e-05, 2.2384e-05, 2.239e-05, 2.2401e-05, 2.2413e-05, 2.2427e-05, 
    2.2439e-05, 2.245e-05, 2.2455e-05, 2.2457e-05, 2.2454e-05, 2.245e-05, 
    2.2445e-05, 2.2443e-05, 2.2443e-05, 2.2446e-05, 2.2454e-05, 2.2464e-05, 
    2.248e-05, 2.2496e-05, 2.2516e-05, 2.2536e-05, 2.2555e-05, 2.2568e-05, 
    2.2577e-05, 2.2563e-05, 2.2543e-05, 2.2517e-05, 2.2495e-05, 2.2474e-05, 
    2.2464e-05, 2.2458e-05, 2.2455e-05, 2.2455e-05, 2.2456e-05, 2.2459e-05, 
    2.2461e-05, 2.2462e-05, 2.2459e-05, 2.2453e-05, 2.2448e-05, 2.2443e-05, 
    2.2438e-05, 2.2435e-05, 2.2432e-05, 2.2429e-05, 2.2424e-05, 2.2416e-05, 
    2.2402e-05, 2.2383e-05, 2.2359e-05, 2.2335e-05, 2.2316e-05, 2.2294e-05, 
    2.2269e-05, 2.2238e-05, 2.2205e-05, 2.2164e-05, 2.213e-05, 2.2102e-05, 
    2.2085e-05, 2.207e-05, 2.206e-05, 2.2047e-05, 2.2031e-05, 2.2009e-05, 
    2.1986e-05, 2.1973e-05, 2.1963e-05, 2.1959e-05, 2.1958e-05, 2.1958e-05, 
    2.1958e-05, 2.1959e-05, 2.196e-05, 2.1957e-05, 2.1952e-05, 2.1937e-05, 
    2.1923e-05, 2.1914e-05, 2.1907e-05, 2.1901e-05, 2.1909e-05, 2.192e-05, 
    2.1935e-05, 2.1944e-05, 2.1951e-05, 2.1951e-05, 2.1948e-05, 2.1943e-05, 
    2.1945e-05, 2.1953e-05, 2.1962e-05, 2.197e-05, 2.1974e-05, 2.1976e-05, 
    2.1975e-05, 2.1992e-05, 2.2018e-05, 2.2073e-05, 2.2142e-05, 2.2225e-05, 
    2.2329e-05, 2.2441e-05, 2.2578e-05, 2.2726e-05, 2.2888e-05, 2.3047e-05, 
    2.3203e-05, 2.3333e-05, 2.3459e-05, 2.3579e-05, 2.37e-05, 2.3819e-05, 
    2.3927e-05, 2.4028e-05, 2.4114e-05, 2.4197e-05, 2.4278e-05, 2.4367e-05, 
    2.4463e-05, 2.4573e-05, 2.4695e-05, 2.4825e-05, 2.496e-05, 2.5091e-05, 
    2.5212e-05, 2.5324e-05, 2.543e-05, 2.5523e-05, 2.562e-05, 2.5737e-05, 
    2.5849e-05, 2.5956e-05, 2.6041e-05, 2.6118e-05, 2.6175e-05, 2.6222e-05, 
    2.6258e-05, 2.6261e-05, 2.6247e-05, 2.6175e-05, 2.6083e-05, 2.5962e-05, 
    2.58e-05, 2.5619e-05, 2.5387e-05, 2.5141e-05, 2.4874e-05, 2.4595e-05, 
    2.4311e-05, 2.4063e-05, 2.3822e-05, 2.3595e-05, 2.3387e-05, 2.3189e-05, 
    2.3004e-05, 2.282e-05, 2.2636e-05, 2.2455e-05, 2.2277e-05, 2.2126e-05, 
    2.1988e-05, 2.1886e-05, 2.1807e-05, 2.1746e-05, 2.1698e-05, 2.1651e-05, 
    2.1599e-05, 2.1542e-05, 2.148e-05, 2.1449e-05, 2.1428e-05, 2.1432e-05, 
    2.1445e-05, 2.1466e-05, 2.1497e-05, 2.153e-05, 2.1565e-05, 2.16e-05, 
    2.1634e-05, 2.1678e-05, 2.1727e-05, 2.179e-05, 2.185e-05, 2.1902e-05, 
    2.1933e-05, 2.1953e-05, 2.1959e-05, 2.1965e-05, 2.1969e-05, 2.1978e-05, 
    2.1988e-05, 2.2003e-05, 2.2017e-05, 2.2027e-05, 2.2032e-05, 2.2035e-05, 
    2.2037e-05, 2.2039e-05, 2.2042e-05, 2.2046e-05, 2.2052e-05, 2.2058e-05, 
    2.2062e-05, 2.2065e-05, 2.2066e-05, 2.2067e-05, 2.2067e-05, 2.2067e-05, 
    2.207e-05, 2.2074e-05, 2.2079e-05, 2.2084e-05, 2.2088e-05, 2.209e-05, 
    2.209e-05, 2.2089e-05, 2.2086e-05, 2.2083e-05, 2.2081e-05, 2.2085e-05, 
    2.2096e-05, 2.2113e-05, 2.2133e-05, 2.2155e-05, 2.2179e-05, 2.2204e-05, 
    2.2232e-05, 2.2262e-05, 2.2299e-05, 2.2336e-05, 2.2369e-05, 2.2393e-05, 
    2.241e-05, 2.2417e-05, 2.2424e-05, 2.2427e-05, 2.2428e-05, 2.2428e-05, 
    2.2428e-05, 2.2427e-05, 2.2427e-05, 2.2426e-05, 2.2426e-05, 2.2427e-05, 
    2.2427e-05, 2.2427e-05, 2.2429e-05, 2.2433e-05, 2.244e-05, 2.2447e-05, 
    2.2454e-05, 2.246e-05, 2.2464e-05, 2.2467e-05, 2.247e-05, 2.2472e-05, 
    2.2474e-05, 2.2477e-05, 2.2475e-05, 2.247e-05, 2.2462e-05, 2.2456e-05, 
    2.2451e-05, 2.2443e-05, 2.2435e-05, 2.2419e-05, 2.2402e-05, 2.2387e-05, 
    2.238e-05, 2.238e-05, 2.2399e-05, 2.2423e-05, 2.2457e-05, 2.2503e-05, 
    2.2559e-05, 2.263e-05, 2.2705e-05, 2.2791e-05, 2.2875e-05, 2.2957e-05, 
    2.3022e-05, 2.3081e-05, 2.3122e-05, 2.3156e-05, 2.3183e-05, 2.3208e-05, 
    2.3232e-05, 2.3253e-05, 2.3272e-05, 2.329e-05, 2.3318e-05, 2.335e-05, 
    2.3391e-05, 2.3434e-05, 2.3478e-05, 2.3504e-05, 2.3524e-05, 2.3524e-05, 
    2.3522e-05, 2.3515e-05, 2.3503e-05, 2.3488e-05, 2.3456e-05, 2.3419e-05, 
    2.3372e-05, 2.3329e-05, 2.3288e-05, 2.3267e-05, 2.3253e-05, 2.3254e-05, 
    2.3258e-05, 2.3264e-05, 2.3259e-05, 2.325e-05, 2.3226e-05, 2.3203e-05, 
    2.318e-05, 2.3162e-05, 2.3147e-05, 2.3141e-05, 2.3138e-05, 2.3138e-05, 
    2.3136e-05, 2.3133e-05, 2.3131e-05, 2.3131e-05, 2.3135e-05, 2.3147e-05, 
    2.3161e-05, 2.3174e-05, 2.3185e-05, 2.3193e-05, 2.3198e-05, 2.3202e-05, 
    2.3206e-05, 2.321e-05, 2.3218e-05, 2.3227e-05, 2.3238e-05, 2.3246e-05, 
    2.3252e-05, 2.3254e-05, 2.3252e-05, 2.3246e-05, 2.323e-05, 2.321e-05, 
    2.3183e-05, 2.315e-05, 2.3114e-05, 2.3085e-05, 2.3061e-05, 2.3051e-05, 
    2.3047e-05, 2.3049e-05, 2.3053e-05, 2.3057e-05, 2.3062e-05, 2.3062e-05, 
    2.306e-05, 2.3044e-05, 2.3024e-05, 2.2989e-05, 2.2956e-05, 2.2924e-05, 
    2.2904e-05, 2.289e-05, 2.2896e-05, 2.2905e-05, 2.2917e-05, 2.2927e-05, 
    2.2937e-05, 2.2945e-05, 2.2953e-05, 2.2961e-05, 2.2972e-05, 2.2983e-05, 
    2.2996e-05, 2.3007e-05, 2.3015e-05, 2.3022e-05, 2.3027e-05, 2.3027e-05, 
    2.3025e-05, 2.302e-05, 2.3012e-05, 2.3002e-05, 2.2991e-05, 2.2981e-05, 
    2.2974e-05, 2.297e-05, 2.2969e-05, 2.2969e-05, 2.2968e-05, 2.2967e-05, 
    2.2963e-05, 2.2957e-05, 2.2945e-05, 2.2931e-05, 2.2909e-05, 2.2885e-05, 
    2.2856e-05, 2.2825e-05, 2.2793e-05, 2.2761e-05, 2.2733e-05, 2.2711e-05, 
    2.2694e-05, 2.2679e-05, 2.267e-05, 2.2662e-05, 2.2658e-05, 2.2659e-05, 
    2.2662e-05, 2.267e-05, 2.2678e-05, 2.2688e-05, 2.2698e-05, 2.2708e-05, 
    2.2716e-05, 2.2723e-05, 2.2723e-05, 2.2721e-05, 2.2716e-05, 2.2709e-05, 
    2.2702e-05, 2.2694e-05, 2.2688e-05, 2.2682e-05, 2.2677e-05, 2.2673e-05, 
    2.267e-05, 2.2668e-05, 2.2667e-05, 2.2667e-05, 2.2667e-05, 2.2667e-05, 
    2.2666e-05, 2.2665e-05, 2.2664e-05, 2.2663e-05, 2.2664e-05, 2.2666e-05, 
    2.2667e-05, 2.2669e-05, 2.2671e-05, 2.2673e-05, 2.2675e-05, 2.2677e-05, 
    2.2679e-05, 2.2681e-05, 2.2686e-05, 2.2694e-05, 2.2706e-05, 2.2719e-05, 
    2.2734e-05, 2.2747e-05, 2.2759e-05, 2.2769e-05, 2.2769e-05, 2.2761e-05, 
    2.2748e-05, 2.2734e-05, 2.2716e-05, 2.2696e-05, 2.2674e-05, 2.2655e-05, 
    2.2638e-05, 2.2624e-05, 2.2611e-05, 2.2598e-05, 2.2588e-05, 2.2579e-05, 
    2.2573e-05, 2.2568e-05, 2.2564e-05, 2.2555e-05, 2.2545e-05, 2.253e-05, 
    2.251e-05, 2.2483e-05, 2.2445e-05, 2.2402e-05, 2.235e-05, 2.2295e-05, 
    2.2231e-05, 2.2159e-05, 2.2082e-05, 2.2011e-05, 2.1944e-05, 2.1887e-05, 
    2.1825e-05, 2.1761e-05, 2.1688e-05, 2.1617e-05, 2.155e-05, 2.1491e-05, 
    2.1436e-05, 2.1379e-05, 2.1318e-05, 2.1243e-05, 2.1153e-05, 2.1049e-05, 
    2.0921e-05, 2.0788e-05, 2.0649e-05, 2.0514e-05, 2.0384e-05, 2.0258e-05, 
    2.0133e-05, 2.0013e-05, 1.9889e-05, 1.9761e-05, 1.9638e-05, 1.9519e-05, 
    1.9427e-05, 1.9339e-05, 1.9259e-05, 1.9178e-05, 1.9096e-05, 1.9025e-05, 
    1.8959e-05, 1.8902e-05, 1.8847e-05, 1.8792e-05, 1.8752e-05, 1.8716e-05, 
    1.8693e-05, 1.8679e-05, 1.8672e-05, 1.8673e-05, 1.8675e-05, 1.8678e-05, 
    1.8685e-05, 1.8694e-05, 1.8707e-05, 1.8722e-05, 1.874e-05, 1.8762e-05, 
    1.8788e-05, 1.8819e-05, 1.8853e-05, 1.8893e-05, 1.893e-05, 1.8964e-05, 
    1.8991e-05, 1.9016e-05, 1.9031e-05, 1.9043e-05, 1.9048e-05, 1.9046e-05, 
    1.9042e-05, 1.903e-05, 1.9019e-05, 1.9008e-05, 1.8998e-05, 1.8988e-05, 
    1.897e-05, 1.8952e-05, 1.8933e-05, 1.8914e-05, 1.8896e-05, 1.8864e-05, 
    1.8825e-05, 1.8772e-05, 1.8725e-05, 1.8681e-05, 1.8668e-05, 1.866e-05, 
    1.8664e-05, 1.8669e-05, 1.8675e-05, 1.8677e-05, 1.8676e-05, 1.8673e-05, 
    1.8674e-05, 1.8678e-05, 1.8687e-05, 1.8697e-05, 1.8704e-05, 1.8711e-05, 
    1.8717e-05, 1.8719e-05, 1.872e-05, 1.8719e-05, 1.872e-05, 1.8723e-05, 
    1.8729e-05, 1.8736e-05, 1.8745e-05, 1.8752e-05, 1.8755e-05, 1.8755e-05, 
    1.8752e-05, 1.8746e-05, 1.8742e-05, 1.8741e-05, 1.8745e-05, 1.8752e-05, 
    1.8765e-05, 1.878e-05, 1.8797e-05, 1.8809e-05, 1.8817e-05, 1.8808e-05, 
    1.8794e-05, 1.8772e-05, 1.8745e-05, 1.8713e-05, 1.8672e-05, 1.8628e-05, 
    1.8577e-05, 1.8529e-05, 1.8484e-05, 1.8459e-05, 1.844e-05, 1.8434e-05, 
    1.843e-05, 1.8431e-05, 1.8436e-05, 1.8441e-05, 1.8448e-05, 1.8454e-05, 
    1.846e-05, 1.8464e-05, 1.8466e-05, 1.8467e-05, 1.8468e-05, 1.8467e-05, 
    1.8462e-05, 1.8456e-05, 1.8448e-05, 1.8439e-05, 1.843e-05, 1.8424e-05, 
    1.842e-05, 1.8416e-05, 1.8412e-05, 1.8409e-05, 1.8407e-05, 1.8404e-05, 
    1.8404e-05, 1.8407e-05, 1.8421e-05, 1.8444e-05, 1.8474e-05, 1.8513e-05, 
    1.8553e-05, 1.8591e-05, 1.8625e-05, 1.8656e-05, 1.8678e-05, 1.8695e-05, 
    1.87e-05, 1.8698e-05, 1.869e-05, 1.8661e-05, 1.8624e-05, 1.8571e-05, 
    1.8512e-05, 1.8446e-05, 1.8384e-05, 1.8325e-05, 1.8282e-05, 1.8244e-05, 
    1.8217e-05, 1.8203e-05, 1.8195e-05, 1.8187e-05, 1.8178e-05, 1.8168e-05, 
    1.8141e-05, 1.8104e-05, 1.8035e-05, 1.7958e-05, 1.7863e-05, 1.776e-05, 
    1.7651e-05, 1.7553e-05, 1.7461e-05, 1.7387e-05, 1.7324e-05, 1.7271e-05, 
    1.7235e-05, 1.7203e-05, 1.7175e-05, 1.7146e-05, 1.7117e-05, 1.709e-05, 
    1.7062e-05, 1.7037e-05, 1.7011e-05, 1.6985e-05, 1.6961e-05, 1.6937e-05, 
    1.6921e-05, 1.6908e-05, 1.6898e-05, 1.6892e-05, 1.6888e-05, 1.6883e-05, 
    1.6877e-05, 1.6867e-05, 1.6855e-05, 1.6841e-05, 1.6824e-05, 1.6807e-05, 
    1.6792e-05, 1.6777e-05, 1.6763e-05, 1.6742e-05, 1.6723e-05, 1.6706e-05, 
    1.6691e-05, 1.6678e-05, 1.667e-05, 1.6663e-05, 1.6657e-05, 1.6649e-05, 
    1.664e-05, 1.6627e-05, 1.6613e-05, 1.6601e-05, 1.6591e-05, 1.6584e-05, 
    1.6582e-05, 1.6583e-05, 1.6589e-05, 1.66e-05, 1.6615e-05, 1.6631e-05, 
    1.6647e-05, 1.6657e-05, 1.6664e-05, 1.6668e-05, 1.6672e-05, 1.6677e-05, 
    1.6683e-05, 1.6687e-05, 1.6688e-05, 1.6687e-05, 1.6683e-05, 1.6674e-05, 
    1.6665e-05, 1.6656e-05, 1.6648e-05, 1.6641e-05, 1.663e-05, 1.6617e-05, 
    1.6597e-05, 1.6579e-05, 1.6562e-05, 1.6548e-05, 1.6535e-05, 1.6522e-05, 
    1.651e-05, 1.6498e-05, 1.6484e-05, 1.647e-05, 1.6457e-05, 1.6446e-05, 
    1.6436e-05, 1.6427e-05, 1.6418e-05, 1.641e-05, 1.6402e-05, 1.6395e-05, 
    1.639e-05, 1.6386e-05, 1.6385e-05, 1.6384e-05, 1.6384e-05, 1.6384e-05, 
    1.6384e-05, 1.6385e-05, 1.6385e-05, 1.6385e-05, 1.6385e-05, 1.6386e-05, 
    1.6387e-05, 1.639e-05, 1.6397e-05, 1.6407e-05, 1.6419e-05, 1.6438e-05, 
    1.646e-05, 1.6488e-05, 1.6525e-05, 1.6567e-05, 1.6621e-05, 1.6677e-05, 
    1.6738e-05, 1.6801e-05, 1.6865e-05, 1.6926e-05, 1.6985e-05, 1.7037e-05, 
    1.708e-05, 1.7117e-05, 1.7144e-05, 1.7167e-05, 1.7184e-05, 1.72e-05, 
    1.7216e-05, 1.723e-05, 1.7244e-05, 1.7254e-05, 1.7263e-05, 1.7269e-05, 
    1.7273e-05, 1.7278e-05, 1.7284e-05, 1.7292e-05, 1.7304e-05, 1.7321e-05, 
    1.7341e-05, 1.7372e-05, 1.7406e-05, 1.7447e-05, 1.7483e-05, 1.7516e-05, 
    1.7532e-05, 1.7543e-05, 1.7543e-05, 1.7542e-05, 1.7541e-05, 1.7556e-05, 
    1.7581e-05, 1.7631e-05, 1.7704e-05, 1.7793e-05, 1.7905e-05, 1.8023e-05, 
    1.8156e-05, 1.8291e-05, 1.8427e-05, 1.856e-05, 1.8692e-05, 1.8826e-05, 
    1.8961e-05, 1.9097e-05, 1.9232e-05, 1.9365e-05, 1.9489e-05, 1.9608e-05, 
    1.972e-05, 1.982e-05, 1.9917e-05, 2.002e-05, 2.0129e-05, 2.0248e-05, 
    2.0385e-05, 2.0528e-05, 2.0678e-05, 2.0829e-05, 2.0983e-05, 2.1146e-05, 
    2.1312e-05, 2.1453e-05, 2.1579e-05, 2.1674e-05, 2.1741e-05, 2.1791e-05, 
    2.1805e-05, 2.1807e-05, 2.1783e-05, 2.174e-05, 2.1682e-05, 2.1605e-05, 
    2.1522e-05, 2.1431e-05, 2.1344e-05, 2.1259e-05, 2.1184e-05, 2.1111e-05, 
    2.1045e-05, 2.0982e-05, 2.0923e-05, 2.0877e-05, 2.0834e-05, 2.0798e-05, 
    2.0767e-05, 2.0742e-05, 2.0724e-05, 2.0709e-05, 2.0696e-05, 2.0681e-05, 
    2.0663e-05, 2.064e-05, 2.0616e-05, 2.0584e-05, 2.055e-05, 2.051e-05, 
    2.0465e-05, 2.0417e-05, 2.0358e-05, 2.0294e-05, 2.0219e-05, 2.014e-05, 
    2.0058e-05, 1.9989e-05, 1.9925e-05, 1.9876e-05, 1.9839e-05, 1.9812e-05, 
    1.9798e-05, 1.9786e-05, 1.9781e-05, 1.9776e-05, 1.9774e-05, 1.9772e-05, 
    1.9771e-05, 1.9769e-05, 1.9767e-05, 1.9763e-05, 1.9755e-05, 1.9746e-05, 
    1.973e-05, 1.9712e-05, 1.969e-05, 1.9665e-05, 1.9638e-05, 1.9607e-05, 
    1.9574e-05, 1.9536e-05, 1.9502e-05, 1.9471e-05, 1.9447e-05, 1.9426e-05, 
    1.9412e-05, 1.9404e-05, 1.9399e-05, 1.9397e-05, 1.9396e-05, 1.9396e-05, 
    1.9392e-05, 1.9386e-05, 1.9375e-05, 1.9363e-05, 1.9351e-05, 1.9339e-05, 
    1.9326e-05, 1.932e-05, 1.9316e-05, 1.9314e-05, 1.9315e-05, 1.9319e-05, 
    1.9326e-05, 1.9335e-05, 1.9345e-05, 1.9356e-05, 1.9368e-05, 1.9382e-05, 
    1.9397e-05, 1.9418e-05, 1.9441e-05, 1.9464e-05, 1.9487e-05, 1.9509e-05, 
    1.9534e-05, 1.9562e-05, 1.9593e-05, 1.9626e-05, 1.966e-05, 1.97e-05, 
    1.9739e-05, 1.9776e-05, 1.9807e-05, 1.9835e-05, 1.9855e-05, 1.9872e-05, 
    1.9885e-05, 1.9897e-05, 1.9908e-05, 1.9919e-05, 1.9928e-05, 1.9936e-05, 
    1.9943e-05, 1.9948e-05, 1.9948e-05, 1.9946e-05, 1.9938e-05, 1.993e-05, 
    1.9921e-05, 1.9912e-05, 1.9906e-05, 1.9911e-05, 1.9922e-05, 1.994e-05, 
    1.9965e-05, 1.9994e-05, 2.0029e-05, 2.0069e-05, 2.0115e-05, 2.017e-05, 
    2.0228e-05, 2.0289e-05, 2.0347e-05, 2.0402e-05, 2.0448e-05, 2.0491e-05, 
    2.0523e-05, 2.0553e-05, 2.0577e-05, 2.0595e-05, 2.061e-05, 2.0618e-05, 
    2.0625e-05, 2.0629e-05, 2.0631e-05, 2.0632e-05, 2.0632e-05, 2.0632e-05, 
    2.0634e-05, 2.0636e-05, 2.064e-05, 2.0645e-05, 2.0651e-05, 2.0657e-05, 
    2.0666e-05, 2.0675e-05, 2.0688e-05, 2.0702e-05, 2.0716e-05, 2.0725e-05, 
    2.0728e-05, 2.0718e-05, 2.0705e-05, 2.0687e-05, 2.0671e-05, 2.0658e-05, 
    2.0654e-05, 2.0654e-05, 2.0661e-05, 2.0667e-05, 2.067e-05, 2.0669e-05, 
    2.0665e-05, 2.0655e-05, 2.0642e-05, 2.0625e-05, 2.0603e-05, 2.0577e-05, 
    2.0542e-05, 2.0505e-05, 2.0462e-05, 2.0414e-05, 2.0363e-05, 2.0311e-05, 
    2.0257e-05, 2.0203e-05, 2.0148e-05, 2.0092e-05, 2.005e-05, 2.0013e-05, 
    1.9987e-05, 1.9967e-05, 1.9951e-05, 1.9943e-05, 1.9937e-05, 1.9934e-05, 
    1.9934e-05, 1.9936e-05, 1.9943e-05, 1.9954e-05, 1.9973e-05, 1.9995e-05, 
    2.0023e-05, 2.0061e-05, 2.0103e-05, 2.0154e-05, 2.0206e-05, 2.0259e-05, 
    2.031e-05, 2.0361e-05, 2.0409e-05, 2.0455e-05, 2.0496e-05, 2.0539e-05, 
    2.0583e-05, 2.0639e-05, 2.0699e-05, 2.0767e-05, 2.0842e-05, 2.0921e-05, 
    2.1013e-05, 2.111e-05, 2.1222e-05, 2.1344e-05, 2.1472e-05, 2.161e-05, 
    2.1751e-05, 2.1904e-05, 2.2056e-05, 2.2209e-05, 2.2338e-05, 2.2458e-05, 
    2.2552e-05, 2.2633e-05, 2.2699e-05, 2.2751e-05, 2.2798e-05, 2.2833e-05, 
    2.2867e-05, 2.2897e-05, 2.2924e-05, 2.2949e-05, 2.2972e-05, 2.2996e-05, 
    2.3019e-05, 2.3044e-05, 2.307e-05, 2.3101e-05, 2.3132e-05, 2.3165e-05, 
    2.3199e-05, 2.3234e-05, 2.3253e-05, 2.3268e-05, 2.3271e-05, 2.3269e-05, 
    2.3264e-05, 2.3259e-05, 2.3257e-05, 2.3261e-05, 2.3273e-05, 2.3293e-05, 
    2.3328e-05, 2.3368e-05, 2.3425e-05, 2.3491e-05, 2.3568e-05, 2.3653e-05, 
    2.3738e-05, 2.382e-05, 2.3895e-05, 2.3966e-05, 2.4027e-05, 2.4086e-05, 
    2.4141e-05, 2.4196e-05, 2.4249e-05, 2.4305e-05, 2.4362e-05, 2.4423e-05, 
    2.4492e-05, 2.4572e-05, 2.4666e-05, 2.4767e-05, 2.4887e-05, 2.5012e-05, 
    2.5146e-05, 2.5283e-05, 2.5421e-05, 2.5546e-05, 2.5664e-05, 2.5767e-05, 
    2.5857e-05, 2.5939e-05, 2.6003e-05, 2.606e-05, 2.6102e-05, 2.6138e-05, 
    2.6168e-05, 2.6192e-05, 2.6213e-05, 2.6229e-05, 2.624e-05, 2.6247e-05, 
    2.6244e-05, 2.6237e-05, 2.622e-05, 2.6201e-05, 2.618e-05, 2.6161e-05, 
    2.6142e-05, 2.6125e-05, 2.6111e-05, 2.6101e-05, 2.6098e-05, 2.6098e-05, 
    2.6108e-05, 2.6119e-05, 2.6131e-05, 2.6139e-05, 2.6144e-05, 2.6145e-05, 
    2.6145e-05, 2.6143e-05, 2.614e-05, 2.6137e-05, 2.6134e-05, 2.6131e-05, 
    2.6126e-05, 2.612e-05, 2.6112e-05, 2.6099e-05, 2.6084e-05, 2.6064e-05, 
    2.6039e-05, 2.6011e-05, 2.5988e-05, 2.5968e-05, 2.5959e-05, 2.5957e-05, 
    2.596e-05, 2.5967e-05, 2.5973e-05, 2.5972e-05, 2.5962e-05, 2.5942e-05, 
    2.5905e-05, 2.5864e-05, 2.5815e-05, 2.5761e-05, 2.5702e-05, 2.5638e-05, 
    2.5573e-05, 2.5513e-05, 2.5455e-05, 2.54e-05, 2.5346e-05, 2.5293e-05, 
    2.5245e-05, 2.5201e-05, 2.5161e-05, 2.5129e-05, 2.51e-05, 2.5081e-05, 
    2.5061e-05, 2.5037e-05, 2.4995e-05, 2.4943e-05, 2.4853e-05, 2.4754e-05, 
    2.4637e-05, 2.4512e-05, 2.4381e-05, 2.4238e-05, 2.4096e-05, 2.3966e-05, 
    2.3854e-05, 2.3757e-05, 2.3693e-05, 2.3641e-05, 2.3621e-05, 2.3612e-05, 
    2.3615e-05, 2.363e-05, 2.3647e-05, 2.3664e-05, 2.3678e-05, 2.3689e-05, 
    2.3695e-05, 2.3698e-05, 2.3696e-05, 2.369e-05, 2.368e-05, 2.3667e-05, 
    2.3653e-05, 2.3635e-05, 2.3617e-05, 2.3597e-05, 2.3578e-05, 2.3558e-05, 
    2.354e-05, 2.3524e-05, 2.3513e-05, 2.3508e-05, 2.3505e-05, 2.3507e-05, 
    2.3509e-05, 2.3512e-05, 2.3514e-05, 2.3516e-05, 2.3519e-05, 2.3524e-05, 
    2.3534e-05, 2.3549e-05, 2.3568e-05, 2.3593e-05, 2.3619e-05, 2.3647e-05, 
    2.3677e-05, 2.3708e-05, 2.3742e-05, 2.3776e-05, 2.3808e-05, 2.3838e-05, 
    2.3865e-05, 2.3885e-05, 2.3902e-05, 2.3914e-05, 2.3923e-05, 2.3931e-05, 
    2.3935e-05, 2.3939e-05, 2.394e-05, 2.3942e-05, 2.3942e-05, 2.3942e-05, 
    2.3942e-05, 2.3943e-05, 2.3943e-05, 2.3944e-05, 2.3945e-05, 2.3945e-05, 
    2.3944e-05, 2.3942e-05, 2.394e-05, 2.3939e-05, 2.3938e-05, 2.3938e-05, 
    2.3938e-05, 2.3938e-05, 2.3938e-05, 2.3938e-05, 2.3937e-05, 2.3935e-05, 
    2.393e-05, 2.3924e-05, 2.3916e-05, 2.3908e-05, 2.3898e-05, 2.3888e-05, 
    2.3878e-05, 2.3868e-05, 2.3856e-05, 2.3843e-05, 2.3826e-05, 2.3809e-05, 
    2.3792e-05, 2.3773e-05, 2.3753e-05, 2.3729e-05, 2.3703e-05, 2.3673e-05, 
    2.364e-05, 2.3606e-05, 2.3573e-05, 2.3539e-05, 2.3507e-05, 2.3473e-05, 
    2.3439e-05, 2.3403e-05, 2.3366e-05, 2.3325e-05, 2.3287e-05, 2.3251e-05, 
    2.322e-05, 2.3191e-05, 2.3167e-05, 2.3145e-05, 2.3125e-05, 2.3106e-05, 
    2.3089e-05, 2.3077e-05, 2.3067e-05, 2.3061e-05, 2.3057e-05, 2.3054e-05, 
    2.3052e-05, 2.3051e-05, 2.305e-05, 2.3048e-05, 2.3044e-05, 2.3038e-05, 
    2.303e-05, 2.3018e-05, 2.3002e-05, 2.2982e-05, 2.2957e-05, 2.293e-05, 
    2.2899e-05, 2.2862e-05, 2.2821e-05, 2.2771e-05, 2.2719e-05, 2.2665e-05, 
    2.2613e-05, 2.2563e-05, 2.2521e-05, 2.2483e-05, 2.2452e-05, 2.2426e-05, 
    2.2403e-05, 2.2385e-05, 2.237e-05, 2.236e-05, 2.2354e-05, 2.2351e-05, 
    2.2351e-05, 2.2351e-05, 2.2353e-05, 2.2354e-05, 2.2354e-05, 2.2352e-05, 
    2.2349e-05, 2.2345e-05, 2.2339e-05, 2.2333e-05, 2.2325e-05, 2.2316e-05, 
    2.2305e-05, 2.2293e-05, 2.2281e-05, 2.2271e-05, 2.2264e-05, 2.2263e-05, 
    2.2265e-05, 2.2271e-05, 2.2278e-05, 2.2286e-05, 2.2296e-05, 2.2306e-05, 
    2.2317e-05, 2.2335e-05, 2.2358e-05, 2.2391e-05, 2.2429e-05, 2.2481e-05, 
    2.2542e-05, 2.2608e-05, 2.2674e-05, 2.2739e-05, 2.2798e-05, 2.2856e-05, 
    2.2914e-05, 2.2967e-05, 2.3019e-05, 2.3063e-05, 2.3104e-05, 2.3141e-05, 
    2.317e-05, 2.3197e-05, 2.3214e-05, 2.3227e-05, 2.3236e-05, 2.3241e-05, 
    2.3244e-05, 2.3244e-05, 2.3244e-05, 2.3244e-05, 2.3243e-05, 2.3243e-05, 
    2.3237e-05, 2.3229e-05, 2.3215e-05, 2.3196e-05, 2.3173e-05, 2.3138e-05, 
    2.31e-05, 2.3055e-05, 2.3008e-05, 2.2959e-05, 2.2909e-05, 2.286e-05, 
    2.2814e-05, 2.2771e-05, 2.273e-05, 2.2688e-05, 2.2644e-05, 2.2592e-05, 
    2.2535e-05, 2.2473e-05, 2.2401e-05, 2.2324e-05, 2.2239e-05, 2.2144e-05, 
    2.2039e-05, 2.1922e-05, 2.1801e-05, 2.1673e-05, 2.1541e-05, 2.1404e-05, 
    2.1269e-05, 2.1137e-05, 2.1037e-05, 2.0952e-05, 2.0891e-05, 2.0855e-05, 
    2.083e-05, 2.083e-05, 2.0836e-05, 2.0853e-05, 2.0876e-05, 2.0901e-05, 
    2.0934e-05, 2.0967e-05, 2.1e-05, 2.1026e-05, 2.1049e-05, 2.1059e-05, 
    2.1064e-05, 2.1058e-05, 2.1045e-05, 2.1028e-05, 2.1002e-05, 2.0978e-05, 
    2.0961e-05, 2.095e-05, 2.0945e-05, 2.0944e-05, 2.0945e-05, 2.0945e-05, 
    2.0941e-05, 2.0932e-05, 2.0911e-05, 2.0884e-05, 2.0841e-05, 2.079e-05, 
    2.0728e-05, 2.065e-05, 2.0568e-05, 2.0476e-05, 2.0388e-05, 2.0306e-05, 
    2.0236e-05, 2.0172e-05, 2.0124e-05, 2.008e-05, 2.0041e-05, 2.0003e-05, 
    1.9967e-05, 1.9925e-05, 1.988e-05, 1.9827e-05, 1.9758e-05, 1.9677e-05, 
    1.9566e-05, 1.9444e-05, 1.9297e-05, 1.9135e-05, 1.8961e-05, 1.8777e-05, 
    1.8594e-05, 1.8422e-05, 1.8264e-05, 1.8117e-05, 1.7993e-05, 1.7876e-05, 
    1.778e-05, 1.7696e-05, 1.7624e-05, 1.7564e-05, 1.7508e-05, 1.7456e-05, 
    1.7405e-05, 1.7357e-05, 1.7312e-05, 1.7267e-05, 1.7229e-05, 1.7194e-05, 
    1.7164e-05, 1.7136e-05, 1.7107e-05, 1.7072e-05, 1.7034e-05, 1.6992e-05, 
    1.6947e-05, 1.6901e-05, 1.685e-05, 1.6798e-05, 1.6742e-05, 1.669e-05, 
    1.6641e-05, 1.6609e-05, 1.6581e-05, 1.6564e-05, 1.6553e-05, 1.6548e-05, 
    1.6551e-05, 1.6555e-05, 1.6562e-05, 1.657e-05, 1.6579e-05, 1.6591e-05, 
    1.6604e-05, 1.662e-05, 1.6641e-05, 1.6666e-05, 1.6699e-05, 1.6736e-05, 
    1.6781e-05, 1.6828e-05, 1.6879e-05, 1.6928e-05, 1.6977e-05, 1.7022e-05, 
    1.7067e-05, 1.7111e-05, 1.715e-05, 1.7186e-05, 1.7204e-05, 1.7215e-05, 
    1.7214e-05, 1.7202e-05, 1.7185e-05, 1.7152e-05, 1.7114e-05, 1.7062e-05, 
    1.6999e-05, 1.6929e-05, 1.6856e-05, 1.6783e-05, 1.6717e-05, 1.6659e-05, 
    1.6606e-05, 1.6568e-05, 1.6535e-05, 1.6517e-05, 1.6508e-05, 1.6509e-05, 
    1.6533e-05, 1.6566e-05, 1.6622e-05, 1.6685e-05, 1.6758e-05, 1.6827e-05, 
    1.689e-05, 1.6925e-05, 1.6949e-05, 1.696e-05, 1.6963e-05, 1.6961e-05, 
    1.6954e-05, 1.6943e-05, 1.6927e-05, 1.6905e-05, 1.6882e-05, 1.6861e-05, 
    1.6844e-05, 1.6834e-05, 1.6831e-05, 1.6833e-05, 1.6844e-05, 1.6856e-05, 
    5.2279e-06, 5.2153e-06, 5.1993e-06, 5.1802e-06, 5.1583e-06, 5.1335e-06, 
    5.1063e-06, 5.0769e-06, 5.0454e-06, 5.0123e-06, 4.9776e-06, 4.9418e-06, 
    4.9049e-06, 4.8673e-06, 4.8293e-06, 4.791e-06, 4.7528e-06, 4.7149e-06, 
    4.6774e-06, 4.6407e-06, 4.605e-06, 4.5704e-06, 4.5371e-06, 4.5054e-06, 
    4.4754e-06, 4.4472e-06, 4.4209e-06, 4.3968e-06, 4.3749e-06, 4.3553e-06, 
    4.3382e-06, 4.3235e-06, 4.3114e-06, 4.302e-06, 4.2954e-06, 4.2916e-06, 
    4.2907e-06, 4.2928e-06, 4.2979e-06, 4.3063e-06, 4.3176e-06, 4.3325e-06, 
    4.3506e-06, 4.3721e-06, 4.3971e-06, 4.4256e-06, 4.4576e-06, 4.493e-06, 
    4.532e-06, 4.5742e-06, 4.6196e-06, 4.668e-06, 4.7191e-06, 4.7725e-06, 
    4.8281e-06, 4.8852e-06, 4.9433e-06, 5.0019e-06, 5.0602e-06, 5.1175e-06, 
    5.1732e-06, 5.2263e-06, 5.2761e-06, 5.3216e-06, 5.3623e-06, 5.3972e-06, 
    5.4259e-06, 5.4475e-06, 5.4617e-06, 5.4681e-06, 5.4663e-06, 5.4564e-06, 
    5.4383e-06, 5.4125e-06, 5.3789e-06, 5.3385e-06, 5.2918e-06, 5.2393e-06, 
    5.1821e-06, 5.1211e-06, 5.0572e-06, 4.9915e-06, 4.9248e-06, 4.8582e-06, 
    4.7926e-06, 4.7289e-06, 4.6679e-06, 4.6103e-06, 4.5567e-06, 4.5076e-06, 
    4.4635e-06, 4.4248e-06, 4.3918e-06, 4.3645e-06, 4.3432e-06, 4.3279e-06, 
    4.3185e-06, 4.315e-06, 4.3171e-06, 4.3247e-06, 4.3375e-06, 4.3552e-06, 
    4.3773e-06, 4.4035e-06, 4.4332e-06, 4.4661e-06, 4.5015e-06, 4.5388e-06, 
    4.5775e-06, 4.6169e-06, 4.6564e-06, 4.6955e-06, 4.7334e-06, 4.7696e-06, 
    4.8035e-06, 4.8346e-06, 4.8624e-06, 4.8866e-06, 4.9069e-06, 4.9229e-06, 
    4.9347e-06, 4.9421e-06, 4.945e-06, 4.9436e-06, 4.9381e-06, 4.9288e-06, 
    4.9158e-06, 4.8996e-06, 4.8806e-06, 4.859e-06, 4.8354e-06, 4.81e-06, 
    4.7834e-06, 4.7557e-06, 4.7275e-06, 4.6988e-06, 4.6701e-06, 4.6413e-06, 
    4.6129e-06, 4.5848e-06, 4.5572e-06, 4.5301e-06, 4.5035e-06, 4.4773e-06, 
    4.4516e-06, 4.4263e-06, 4.4015e-06, 4.3771e-06, 4.3529e-06, 4.329e-06, 
    4.3055e-06, 4.2823e-06, 4.2595e-06, 4.2371e-06, 4.2151e-06, 4.1936e-06, 
    4.1728e-06, 4.1527e-06, 4.1334e-06, 4.1149e-06, 4.0973e-06, 4.0807e-06, 
    4.0652e-06, 4.0508e-06, 4.0375e-06, 4.0253e-06, 4.0142e-06, 4.0043e-06, 
    3.9954e-06, 3.9877e-06, 3.9809e-06, 3.975e-06, 3.9701e-06, 3.966e-06, 
    3.9626e-06, 3.9599e-06, 3.9578e-06, 3.9562e-06, 3.955e-06, 3.9543e-06, 
    3.9538e-06, 3.9535e-06, 3.9534e-06, 3.9534e-06, 3.9533e-06, 3.9533e-06, 
    3.953e-06, 3.9525e-06, 3.9515e-06, 3.9501e-06, 3.9482e-06, 3.9454e-06, 
    3.9418e-06, 3.9371e-06, 3.9315e-06, 3.9245e-06, 3.9163e-06, 3.9067e-06, 
    3.8957e-06, 3.8833e-06, 3.8694e-06, 3.8542e-06, 3.8376e-06, 3.8198e-06, 
    3.801e-06, 3.7812e-06, 3.7605e-06, 3.7392e-06, 3.7173e-06, 3.6949e-06, 
    3.6724e-06, 3.6496e-06, 3.6267e-06, 3.6038e-06, 3.581e-06, 3.5583e-06, 
    3.5357e-06, 3.5134e-06, 3.4914e-06, 3.4697e-06, 3.4483e-06, 3.4274e-06, 
    3.407e-06, 3.3872e-06, 3.3681e-06, 3.3498e-06, 3.3324e-06, 3.3161e-06, 
    3.3009e-06, 3.287e-06, 3.2745e-06, 3.2635e-06, 3.2541e-06, 3.2465e-06, 
    3.2406e-06, 3.2365e-06, 3.2343e-06, 3.234e-06, 3.2356e-06, 3.2391e-06, 
    3.2445e-06, 3.2516e-06, 3.2605e-06, 3.2711e-06, 3.2831e-06, 3.2966e-06, 
    3.3115e-06, 3.3275e-06, 3.3446e-06, 3.3626e-06, 3.3814e-06, 3.4008e-06, 
    3.4208e-06, 3.4413e-06, 3.4621e-06, 3.4832e-06, 3.5046e-06, 3.5262e-06, 
    3.548e-06, 3.57e-06, 3.5922e-06, 3.6147e-06, 3.6374e-06, 3.6604e-06, 
    3.6837e-06, 3.7074e-06, 3.7313e-06, 3.7556e-06, 3.78e-06, 3.8046e-06, 
    3.8292e-06, 3.8536e-06, 3.8776e-06, 3.901e-06, 3.9236e-06, 3.945e-06, 
    3.9648e-06, 3.983e-06, 3.9989e-06, 4.0126e-06, 4.0234e-06, 4.0314e-06, 
    4.0361e-06, 4.0374e-06, 4.0353e-06, 4.0296e-06, 4.0204e-06, 4.0077e-06, 
    3.9917e-06, 3.9725e-06, 3.9504e-06, 3.9257e-06, 3.8987e-06, 3.8698e-06, 
    3.8393e-06, 3.8077e-06, 3.775e-06, 3.742e-06, 3.7086e-06, 3.6754e-06, 
    3.6425e-06, 3.6101e-06, 3.5783e-06, 3.5474e-06, 3.5174e-06, 3.4883e-06, 
    3.4602e-06, 3.4331e-06, 3.4069e-06, 3.3816e-06, 3.3574e-06, 3.3339e-06, 
    3.3113e-06, 3.2896e-06, 3.2685e-06, 3.2483e-06, 3.2287e-06, 3.2099e-06, 
    3.1918e-06, 3.1743e-06, 3.1577e-06, 3.1416e-06, 3.1263e-06, 3.1117e-06, 
    3.0978e-06, 3.0846e-06, 3.0721e-06, 3.0604e-06, 3.0494e-06, 3.0391e-06, 
    3.0295e-06, 3.0208e-06, 3.0129e-06, 3.0058e-06, 2.9996e-06, 2.9943e-06, 
    2.9899e-06, 2.9865e-06, 2.9841e-06, 2.9827e-06, 2.9823e-06, 2.9828e-06, 
    2.9843e-06, 2.9868e-06, 2.9901e-06, 2.9943e-06, 2.9992e-06, 3.0049e-06, 
    3.0111e-06, 3.0178e-06, 3.025e-06, 3.0325e-06, 3.0403e-06, 3.0483e-06, 
    3.0565e-06, 3.0647e-06, 3.0729e-06, 3.0812e-06, 3.0893e-06, 3.0973e-06, 
    3.1053e-06, 3.1131e-06, 3.1207e-06, 3.1283e-06, 3.1356e-06, 3.1428e-06, 
    3.1499e-06, 3.1568e-06, 3.1636e-06, 3.1703e-06, 3.1769e-06, 3.1835e-06, 
    3.1902e-06, 3.1969e-06, 3.2038e-06, 3.2108e-06, 3.2181e-06, 3.2257e-06, 
    3.2337e-06, 3.2421e-06, 3.251e-06, 3.2604e-06, 3.2703e-06, 3.2806e-06, 
    3.2914e-06, 3.3025e-06, 3.3139e-06, 3.3255e-06, 3.3371e-06, 3.3485e-06, 
    3.3595e-06, 3.3699e-06, 3.3795e-06, 3.3879e-06, 3.3951e-06, 3.4006e-06, 
    3.4044e-06, 3.4062e-06, 3.4058e-06, 3.4031e-06, 3.398e-06, 3.3904e-06, 
    3.3805e-06, 3.3682e-06, 3.3536e-06, 3.3369e-06, 3.3184e-06, 3.2981e-06, 
    3.2765e-06, 3.2537e-06, 3.2301e-06, 3.206e-06, 3.1816e-06, 3.1573e-06, 
    3.1333e-06, 3.1098e-06, 3.087e-06, 3.0652e-06, 3.0446e-06, 3.0252e-06, 
    3.0071e-06, 2.9904e-06, 2.9752e-06, 2.9614e-06, 2.949e-06, 2.9381e-06, 
    2.9284e-06, 2.9201e-06, 2.9129e-06, 2.9067e-06, 2.9015e-06, 2.8971e-06, 
    2.8934e-06, 2.8902e-06, 2.8875e-06, 2.8851e-06, 2.883e-06, 2.8809e-06, 
    2.879e-06, 2.877e-06, 2.8749e-06, 2.8728e-06, 2.8706e-06, 2.8682e-06, 
    2.8658e-06, 2.8634e-06, 2.8611e-06, 2.8587e-06, 2.8565e-06, 2.8545e-06, 
    2.8527e-06, 2.8513e-06, 2.8501e-06, 2.8492e-06, 2.8486e-06, 2.8483e-06, 
    2.8482e-06, 2.8483e-06, 2.8483e-06, 2.8483e-06, 2.8482e-06, 2.8476e-06, 
    2.8466e-06, 2.845e-06, 2.8427e-06, 2.8395e-06, 2.8353e-06, 2.83e-06, 
    2.8237e-06, 2.8162e-06, 2.8076e-06, 2.798e-06, 2.7874e-06, 2.7759e-06, 
    2.7639e-06, 2.7512e-06, 2.7383e-06, 2.7254e-06, 2.7125e-06, 2.7001e-06, 
    2.6883e-06, 2.6774e-06, 2.6676e-06, 2.659e-06, 2.6519e-06, 2.6464e-06, 
    2.6426e-06, 2.6406e-06, 2.6405e-06, 2.6423e-06, 2.646e-06, 2.6515e-06, 
    2.6588e-06, 2.6678e-06, 2.6782e-06, 2.6898e-06, 2.7026e-06, 2.7162e-06, 
    2.7303e-06, 2.7447e-06, 2.7591e-06, 2.773e-06, 2.7864e-06, 2.7988e-06, 
    2.81e-06, 2.8198e-06, 2.8279e-06, 2.8341e-06, 2.8384e-06, 2.8407e-06, 
    2.841e-06, 2.839e-06, 2.8351e-06, 2.8293e-06, 2.8216e-06, 2.8121e-06, 
    2.8012e-06, 2.7888e-06, 2.7751e-06, 2.7604e-06, 2.7448e-06, 2.7285e-06, 
    2.7115e-06, 2.6942e-06, 2.6765e-06, 2.6587e-06, 2.6408e-06, 2.623e-06, 
    2.6055e-06, 2.5882e-06, 2.5714e-06, 2.5552e-06, 2.5395e-06, 2.5247e-06, 
    2.5107e-06, 2.4976e-06, 2.4856e-06, 2.4748e-06, 2.4651e-06, 2.4567e-06, 
    2.4496e-06, 2.4438e-06, 2.4394e-06, 2.4364e-06, 2.4346e-06, 2.4342e-06, 
    2.435e-06, 2.437e-06, 2.4399e-06, 2.4439e-06, 2.4487e-06, 2.4542e-06, 
    2.4602e-06, 2.4667e-06, 2.4735e-06, 2.4804e-06, 2.4875e-06, 2.4946e-06, 
    2.5017e-06, 2.5086e-06, 2.5153e-06, 2.522e-06, 2.5285e-06, 2.5348e-06, 
    2.5412e-06, 2.5475e-06, 2.5539e-06, 2.5605e-06, 2.5673e-06, 2.5743e-06, 
    2.5816e-06, 2.5892e-06, 2.5971e-06, 2.6054e-06, 2.6139e-06, 2.6226e-06, 
    2.6313e-06, 2.64e-06, 2.6486e-06, 2.6568e-06, 2.6644e-06, 2.6714e-06, 
    2.6774e-06, 2.6823e-06, 2.6858e-06, 2.6878e-06, 2.6881e-06, 2.6865e-06, 
    2.683e-06, 2.6775e-06, 2.6699e-06, 2.6602e-06, 2.6486e-06, 2.6351e-06, 
    2.6199e-06, 2.603e-06, 2.5849e-06, 2.5658e-06, 2.5458e-06, 2.5254e-06, 
    2.5049e-06, 2.4844e-06, 2.4644e-06, 2.445e-06, 2.4266e-06, 2.4094e-06, 
    2.3936e-06, 2.3792e-06, 2.3665e-06, 2.3556e-06, 2.3464e-06, 2.339e-06, 
    2.3333e-06, 2.3294e-06, 2.327e-06, 2.3262e-06, 2.3266e-06, 2.3283e-06, 
    2.3311e-06, 2.3346e-06, 2.3387e-06, 2.3433e-06, 2.348e-06, 2.3528e-06, 
    2.3575e-06, 2.3618e-06, 2.3657e-06, 2.369e-06, 2.3716e-06, 2.3734e-06, 
    2.3745e-06, 2.3749e-06, 2.3744e-06, 2.3733e-06, 2.3715e-06, 2.3692e-06, 
    2.3664e-06, 2.3633e-06, 2.3599e-06, 2.3565e-06, 2.3531e-06, 2.3498e-06, 
    2.3468e-06, 2.3443e-06, 2.3422e-06, 2.3406e-06, 2.3397e-06, 2.3395e-06, 
    2.34e-06, 2.3412e-06, 2.3433e-06, 2.346e-06, 2.3496e-06, 2.3538e-06, 
    2.3586e-06, 2.3641e-06, 2.37e-06, 2.3764e-06, 2.3831e-06, 2.39e-06, 
    2.3971e-06, 2.4041e-06, 2.411e-06, 2.4176e-06, 2.4239e-06, 2.4297e-06, 
    2.4349e-06, 2.4394e-06, 2.4431e-06, 2.446e-06, 2.448e-06, 2.449e-06, 
    2.449e-06, 2.448e-06, 2.4459e-06, 2.4428e-06, 2.4388e-06, 2.4337e-06, 
    2.4277e-06, 2.4208e-06, 2.413e-06, 2.4044e-06, 2.3949e-06, 2.3848e-06, 
    2.3739e-06, 2.3624e-06, 2.3504e-06, 2.3379e-06, 2.3249e-06, 2.3115e-06, 
    2.2979e-06, 2.284e-06, 2.2701e-06, 2.2562e-06, 2.2424e-06, 2.2288e-06, 
    2.2155e-06, 2.2027e-06, 2.1903e-06, 2.1787e-06, 2.1677e-06, 2.1576e-06, 
    2.1485e-06, 2.1404e-06, 2.1333e-06, 2.1274e-06, 2.1227e-06, 2.1191e-06, 
    2.1168e-06, 2.1158e-06, 2.1159e-06, 2.1172e-06, 2.1197e-06, 2.1232e-06, 
    2.1276e-06, 2.133e-06, 2.1392e-06, 2.1459e-06, 2.1532e-06, 2.161e-06, 
    2.1689e-06, 2.1769e-06, 2.1848e-06, 2.1926e-06, 2.2e-06, 2.207e-06, 
    2.2134e-06, 2.2192e-06, 2.2244e-06, 2.2288e-06, 2.2325e-06, 2.2354e-06, 
    2.2377e-06, 2.2393e-06, 2.2403e-06, 2.2406e-06, 2.2405e-06, 2.2399e-06, 
    2.2389e-06, 2.2375e-06, 2.2358e-06, 2.2338e-06, 2.2316e-06, 2.2292e-06, 
    2.2265e-06, 2.2238e-06, 2.2209e-06, 2.2178e-06, 2.2146e-06, 2.2114e-06, 
    2.2081e-06, 2.2049e-06, 2.2017e-06, 2.1986e-06, 2.1957e-06, 2.1931e-06, 
    2.1908e-06, 2.1888e-06, 2.1873e-06, 2.1862e-06, 2.1857e-06, 2.1858e-06, 
    2.1864e-06, 2.1877e-06, 2.1895e-06, 2.1918e-06, 2.1947e-06, 2.198e-06, 
    2.2017e-06, 2.2057e-06, 2.2098e-06, 2.214e-06, 2.2181e-06, 2.222e-06, 
    2.2256e-06, 2.2287e-06, 2.2311e-06, 2.2329e-06, 2.2338e-06, 2.2339e-06, 
    2.233e-06, 2.2311e-06, 2.2281e-06, 2.2242e-06, 2.2192e-06, 2.2134e-06, 
    2.2067e-06, 2.1993e-06, 2.1912e-06, 2.1826e-06, 2.1736e-06, 2.1644e-06, 
    2.155e-06, 2.1457e-06, 2.1365e-06, 2.1275e-06, 2.119e-06, 2.111e-06, 
    2.1035e-06, 2.0966e-06, 2.0905e-06, 2.0851e-06, 2.0804e-06, 2.0766e-06, 
    2.0735e-06, 2.0713e-06, 2.0697e-06, 2.0688e-06, 2.0686e-06, 2.0689e-06, 
    2.0697e-06, 2.0709e-06, 2.0724e-06, 2.0741e-06, 2.0759e-06, 2.0778e-06, 
    2.0796e-06, 2.0813e-06, 2.0827e-06, 2.0839e-06, 2.0848e-06, 2.0853e-06, 
    2.0855e-06, 2.0853e-06, 2.0848e-06, 2.0839e-06, 2.0828e-06, 2.0814e-06, 
    2.0798e-06, 2.0781e-06, 2.0762e-06, 2.0743e-06, 2.0725e-06, 2.0706e-06, 
    2.0688e-06, 2.0671e-06, 2.0655e-06, 2.0641e-06, 2.0627e-06, 2.0615e-06, 
    2.0604e-06, 2.0594e-06, 2.0585e-06, 2.0576e-06, 2.0569e-06, 2.0562e-06, 
    2.0555e-06, 2.0548e-06, 2.0542e-06, 2.0537e-06, 2.0531e-06, 2.0526e-06, 
    2.0521e-06, 2.0516e-06, 2.0512e-06, 2.0508e-06, 2.0504e-06, 2.05e-06, 
    2.0497e-06, 2.0493e-06, 2.0489e-06, 2.0486e-06, 2.0481e-06, 2.0477e-06, 
    2.0471e-06, 2.0465e-06, 2.0458e-06, 2.045e-06, 2.0441e-06, 2.0431e-06, 
    2.0421e-06, 2.0409e-06, 2.0396e-06, 2.0383e-06, 2.0369e-06, 2.0355e-06, 
    2.0341e-06, 2.0326e-06, 2.0312e-06, 2.0298e-06, 2.0284e-06, 2.027e-06, 
    2.0257e-06, 2.0245e-06, 2.0233e-06, 2.0222e-06, 2.0211e-06, 2.0202e-06, 
    2.0193e-06, 2.0185e-06, 2.0178e-06, 2.0172e-06, 2.0168e-06, 2.0165e-06, 
    2.0163e-06, 2.0164e-06, 2.0166e-06, 2.017e-06, 2.0177e-06, 2.0186e-06, 
    2.0198e-06, 2.0212e-06, 2.0229e-06, 2.0248e-06, 2.0269e-06, 2.0292e-06, 
    2.0317e-06, 2.0343e-06, 2.037e-06, 2.0397e-06, 2.0423e-06, 2.0449e-06, 
    2.0474e-06, 2.0496e-06, 2.0516e-06, 2.0533e-06, 2.0546e-06, 2.0555e-06, 
    2.0561e-06, 2.0562e-06, 2.0559e-06, 2.0552e-06, 2.0542e-06, 2.0527e-06, 
    2.0509e-06, 2.0488e-06, 2.0465e-06, 2.044e-06, 2.0414e-06, 2.0386e-06, 
    2.036e-06, 2.0333e-06, 2.0308e-06, 2.0284e-06, 2.0262e-06, 2.0242e-06, 
    2.0225e-06, 2.0211e-06, 2.0199e-06, 2.019e-06, 2.0185e-06, 2.0182e-06, 
    2.0181e-06, 2.0183e-06, 2.0187e-06, 2.0192e-06, 2.0199e-06, 2.0207e-06, 
    2.0215e-06, 2.0224e-06, 2.0233e-06, 2.0241e-06, 2.025e-06, 2.0257e-06, 
    2.0264e-06, 2.0271e-06, 2.0276e-06, 2.0281e-06, 2.0285e-06, 2.0289e-06, 
    2.0292e-06, 2.0295e-06, 2.0297e-06, 2.0299e-06, 2.0301e-06, 2.0303e-06, 
    2.0304e-06, 2.0305e-06, 2.0306e-06, 2.0306e-06, 2.0306e-06, 2.0305e-06, 
    2.0304e-06, 2.0302e-06, 2.0299e-06, 2.0295e-06, 2.029e-06, 2.0284e-06, 
    2.0277e-06, 2.0269e-06, 2.026e-06, 2.0251e-06, 2.0241e-06, 2.0229e-06, 
    2.0218e-06, 2.0207e-06, 2.0195e-06, 2.0183e-06, 2.0171e-06, 2.0159e-06, 
    2.0147e-06, 2.0136e-06, 2.0124e-06, 2.0113e-06, 2.0102e-06, 2.009e-06, 
    2.0079e-06, 2.0068e-06, 2.0056e-06, 2.0045e-06, 2.0032e-06, 2.002e-06, 
    2.0006e-06, 1.9992e-06, 1.9977e-06, 1.9962e-06, 1.9945e-06, 1.9928e-06, 
    1.991e-06, 1.989e-06, 1.987e-06, 1.9849e-06, 1.9826e-06, 1.9803e-06, 
    1.9779e-06, 1.9754e-06, 1.9728e-06, 1.9701e-06, 1.9675e-06, 1.9647e-06, 
    1.962e-06, 1.9593e-06, 1.9567e-06, 1.9541e-06, 1.9517e-06, 1.9494e-06, 
    1.9472e-06, 1.9453e-06, 1.9436e-06, 1.9421e-06, 1.9409e-06, 1.94e-06, 
    1.9393e-06, 1.939e-06, 1.939e-06, 1.9393e-06, 1.9399e-06, 1.9408e-06, 
    1.9419e-06, 1.9433e-06, 1.9448e-06, 1.9466e-06, 1.9484e-06, 1.9504e-06, 
    1.9525e-06, 1.9547e-06, 1.9569e-06, 1.9591e-06, 1.9612e-06, 1.9634e-06, 
    1.9654e-06, 1.9674e-06, 1.9693e-06, 1.9712e-06, 1.9729e-06, 1.9745e-06, 
    1.9759e-06, 1.9773e-06, 1.9785e-06, 1.9796e-06, 1.9806e-06, 1.9815e-06, 
    1.9823e-06, 1.9829e-06, 1.9834e-06, 1.9839e-06, 1.9842e-06, 1.9844e-06, 
    1.9846e-06, 1.9846e-06, 1.9846e-06, 1.9844e-06, 1.9843e-06, 1.984e-06, 
    1.9837e-06, 1.9833e-06, 1.9828e-06, 1.9823e-06, 1.9818e-06, 1.9812e-06, 
    1.9806e-06, 1.9799e-06, 1.9792e-06, 1.9784e-06, 1.9776e-06, 1.9768e-06, 
    1.9759e-06, 1.975e-06, 1.974e-06, 1.973e-06, 1.9719e-06, 1.9708e-06, 
    1.9696e-06, 1.9683e-06, 1.967e-06, 1.9656e-06, 1.9641e-06, 1.9625e-06, 
    1.9609e-06, 1.9592e-06, 1.9575e-06, 1.9558e-06, 1.954e-06, 1.9523e-06, 
    1.9506e-06, 1.9488e-06, 1.9472e-06, 1.9456e-06, 1.944e-06, 1.9426e-06, 
    1.9412e-06, 1.94e-06, 1.9389e-06, 1.9378e-06, 1.9369e-06, 1.9361e-06, 
    1.9355e-06, 1.9349e-06, 1.9344e-06, 1.9341e-06, 1.9339e-06, 1.9338e-06, 
    1.9338e-06, 1.9339e-06, 1.9341e-06, 1.9344e-06, 1.9349e-06, 1.9354e-06, 
    1.9361e-06, 1.9369e-06, 1.9377e-06, 1.9387e-06, 1.9396e-06, 1.9407e-06, 
    1.9419e-06, 1.943e-06, 1.9441e-06, 1.9452e-06, 1.9463e-06, 1.9473e-06, 
    1.9482e-06, 1.949e-06, 1.9496e-06, 1.95e-06, 1.9503e-06, 1.9504e-06, 
    1.9503e-06, 1.95e-06, 1.9496e-06, 1.9489e-06, 1.9481e-06, 1.9472e-06, 
    1.9461e-06, 1.945e-06, 1.9438e-06, 1.9425e-06, 1.9413e-06, 1.94e-06, 
    1.9389e-06, 1.9377e-06, 1.9367e-06, 1.9358e-06, 1.9349e-06, 1.9342e-06, 
    1.9336e-06, 1.9332e-06, 1.9329e-06, 1.9326e-06, 1.9325e-06, 1.9325e-06, 
    1.9326e-06, 1.9328e-06, 1.933e-06, 1.9332e-06, 1.9336e-06, 1.9339e-06, 
    1.9343e-06, 1.9347e-06, 1.9351e-06, 1.9354e-06, 1.9358e-06, 1.9362e-06, 
    1.9365e-06, 1.9369e-06, 1.9372e-06, 1.9375e-06, 1.9378e-06, 1.938e-06, 
    1.9382e-06, 1.9382e-06, 1.9383e-06, 1.9383e-06, 1.9381e-06, 1.9379e-06, 
    1.9376e-06, 1.9371e-06, 1.9365e-06, 1.9357e-06, 1.9348e-06, 1.9338e-06, 
    1.9326e-06, 1.9314e-06, 1.9301e-06, 1.9288e-06, 1.9275e-06, 1.9263e-06, 
    1.9253e-06, 1.9244e-06, 1.9239e-06, 1.9236e-06, 1.9238e-06, 1.9244e-06, 
    1.9255e-06, 1.9271e-06, 1.9292e-06, 1.9319e-06, 1.9351e-06, 1.9388e-06, 
    1.943e-06, 1.9475e-06, 1.9523e-06, 1.9573e-06, 1.9623e-06, 1.9673e-06, 
    1.9721e-06, 1.9765e-06, 1.9805e-06, 1.9839e-06, 1.9867e-06, 1.9886e-06, 
    1.9897e-06, 1.99e-06, 1.9893e-06, 1.9877e-06, 1.9853e-06, 1.982e-06, 
    1.978e-06, 1.9734e-06, 1.9682e-06, 1.9625e-06, 1.9566e-06, 1.9505e-06, 
    1.9443e-06, 1.9382e-06, 1.9323e-06, 1.9266e-06, 1.9212e-06, 1.9163e-06, 
    1.9118e-06, 1.9078e-06, 1.9043e-06, 1.9014e-06, 1.899e-06, 1.8972e-06, 
    1.8959e-06, 1.8951e-06, 1.8948e-06, 1.8949e-06, 1.8955e-06, 1.8964e-06, 
    1.8978e-06, 1.8995e-06, 1.9014e-06, 1.9037e-06, 1.9062e-06, 1.9089e-06, 
    1.9118e-06, 1.9149e-06, 1.9181e-06, 1.9214e-06, 1.9248e-06, 1.9282e-06, 
    1.9317e-06, 1.9352e-06, 1.9386e-06, 1.942e-06, 1.9452e-06, 1.9484e-06, 
    1.9514e-06, 1.9542e-06, 1.9569e-06, 1.9593e-06, 1.9616e-06, 1.9635e-06, 
    1.9653e-06, 1.9667e-06, 1.9679e-06, 1.9688e-06, 1.9695e-06, 1.9699e-06, 
    1.97e-06, 1.9699e-06, 1.9695e-06, 1.9689e-06, 1.9681e-06, 1.9671e-06, 
    1.9659e-06, 1.9645e-06, 1.9629e-06, 1.9612e-06, 1.9593e-06, 1.9573e-06, 
    1.9552e-06, 1.9528e-06, 1.9504e-06, 1.9479e-06, 1.9453e-06, 1.9425e-06, 
    1.9397e-06, 1.9368e-06, 1.9338e-06, 1.9307e-06, 1.9275e-06, 1.9242e-06, 
    1.9209e-06, 1.9176e-06, 1.9141e-06, 1.9107e-06, 1.9071e-06, 1.9036e-06, 
    1.9001e-06, 1.8966e-06, 1.8932e-06, 1.8898e-06, 1.8865e-06, 1.8834e-06, 
    1.8804e-06, 1.8775e-06, 1.8749e-06, 1.8725e-06, 1.8704e-06, 1.8685e-06, 
    1.8669e-06, 1.8656e-06, 1.8646e-06, 1.8638e-06, 1.8634e-06, 1.8633e-06, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_opt_sigma =
  0.00134, 0.0013437, 0.0013472, 0.0013502, 0.0013528, 0.0013553, 0.0013573, 
    0.0013592, 0.0013606, 0.0013618, 0.0013628, 0.0013638, 0.0013647, 
    0.0013655, 0.0013662, 0.0013668, 0.0013673, 0.0013676, 0.0013676, 
    0.0013673, 0.0013668, 0.001366, 0.0013652, 0.0013643, 0.0013634, 
    0.0013624, 0.0013616, 0.0013608, 0.0013603, 0.0013599, 0.0013597, 
    0.0013598, 0.0013601, 0.0013607, 0.0013615, 0.0013625, 0.0013636, 
    0.0013649, 0.0013663, 0.0013677, 0.0013691, 0.0013704, 0.0013716, 
    0.0013726, 0.0013735, 0.0013743, 0.0013749, 0.0013755, 0.001376, 
    0.0013765, 0.001377, 0.0013775, 0.0013781, 0.0013786, 0.0013792, 
    0.0013798, 0.0013805, 0.0013811, 0.0013818, 0.0013824, 0.0013831, 
    0.0013838, 0.0013845, 0.001385, 0.0013855, 0.001386, 0.0013865, 
    0.0013871, 0.0013877, 0.0013883, 0.001389, 0.0013898, 0.0013906, 
    0.0013915, 0.0013924, 0.0013933, 0.0013942, 0.001395, 0.0013956, 
    0.001396, 0.001396, 0.0013959, 0.0013956, 0.0013953, 0.0013949, 
    0.0013946, 0.0013943, 0.0013939, 0.0013934, 0.0013928, 0.0013922, 
    0.0013916, 0.0013911, 0.0013906, 0.0013902, 0.0013896, 0.0013891, 
    0.0013884, 0.0013878, 0.0013871, 0.0013865, 0.001386, 0.0013857, 
    0.0013854, 0.0013852, 0.0013851, 0.001385, 0.0013851, 0.0013852, 
    0.0013853, 0.0013852, 0.0013852, 0.0013849, 0.0013846, 0.0013842, 
    0.0013837, 0.0013832, 0.0013827, 0.0013821, 0.0013816, 0.0013811, 
    0.0013807, 0.0013804, 0.0013801, 0.0013799, 0.0013797, 0.0013796, 
    0.0013795, 0.0013795, 0.0013795, 0.0013795, 0.0013795, 0.0013796, 
    0.0013796, 0.0013797, 0.0013798, 0.0013799, 0.00138, 0.0013802, 
    0.0013803, 0.0013804, 0.0013804, 0.0013803, 0.0013802, 0.0013798, 
    0.0013792, 0.0013784, 0.0013771, 0.0013757, 0.001374, 0.0013722, 
    0.0013705, 0.0013691, 0.0013679, 0.0013671, 0.0013666, 0.0013664, 
    0.0013664, 0.0013667, 0.0013671, 0.0013675, 0.0013677, 0.0013677, 
    0.0013675, 0.0013665, 0.0013653, 0.001363, 0.00136, 0.0013562, 0.0013509, 
    0.0013451, 0.0013377, 0.0013293, 0.0013198, 0.0013088, 0.0012971, 
    0.001284, 0.0012702, 0.0012555, 0.0012398, 0.0012235, 0.0012061, 
    0.0011881, 0.0011692, 0.0011493, 0.0011287, 0.0011067, 0.0010843, 
    0.0010614, 0.0010386, 0.0010157, 0.0009934, 0.00097129, 0.00095024, 
    0.00093045, 0.0009114, 0.00089528, 0.00088002, 0.00086727, 0.0008562, 
    0.00084648, 0.00083964, 0.00083371, 0.00082995, 0.00082722, 0.00082546, 
    0.00082474, 0.00082431, 0.00082429, 0.00082424, 0.00082417, 0.00082376, 
    0.00082321, 0.00082216, 0.00082093, 0.00081946, 0.00081761, 0.0008156, 
    0.00081304, 0.00081032, 0.00080734, 0.00080406, 0.00080064, 0.00079656, 
    0.00079224, 0.00078745, 0.0007822, 0.00077669, 0.0007708, 0.00076483, 
    0.00075876, 0.00075272, 0.0007467, 0.00074081, 0.00073502, 0.00072958, 
    0.00072453, 0.00071978, 0.00071565, 0.0007117, 0.00070818, 0.00070493, 
    0.00070195, 0.00069941, 0.00069702, 0.00069506, 0.00069329, 0.00069174, 
    0.00069044, 0.00068923, 0.00068813, 0.00068708, 0.00068611, 0.00068523, 
    0.00068439, 0.00068375, 0.00068319, 0.00068276, 0.00068241, 0.00068211, 
    0.00068191, 0.00068175, 0.00068167, 0.00068165, 0.00068165, 0.00068167, 
    0.00068169, 0.00068171, 0.00068173, 0.00068175, 0.00068176, 0.00068177, 
    0.00068176, 0.00068176, 0.00068177, 0.00068179, 0.0006818, 0.00068183, 
    0.00068185, 0.00068187, 0.0006819, 0.00068192, 0.00068193, 0.00068194, 
    0.00068194, 0.00068194, 0.00068192, 0.0006819, 0.00068186, 0.00068182, 
    0.00068175, 0.00068168, 0.00068161, 0.00068153, 0.00068144, 0.00068136, 
    0.00068128, 0.0006812, 0.00068112, 0.00068106, 0.00068101, 0.00068096, 
    0.00068093, 0.00068091, 0.00068089, 0.00068087, 0.00068087, 0.00068088, 
    0.00068089, 0.0006809, 0.00068091, 0.00068091, 0.00068091, 0.0006809, 
    0.00068088, 0.00068084, 0.0006808, 0.00068074, 0.00068067, 0.0006806, 
    0.00068052, 0.00068044, 0.00068036, 0.00068027, 0.00068018, 0.00068009, 
    0.00067999, 0.00067988, 0.00067978, 0.00067966, 0.00067953, 0.00067939, 
    0.00067923, 0.00067907, 0.0006789, 0.00067872, 0.00067852, 0.00067833, 
    0.00067814, 0.00067796, 0.00067778, 0.00067762, 0.00067746, 0.00067731, 
    0.0006772, 0.00067711, 0.00067706, 0.00067703, 0.00067701, 0.00067702, 
    0.00067704, 0.00067707, 0.00067709, 0.0006771, 0.00067708, 0.00067704, 
    0.00067695, 0.00067682, 0.00067664, 0.00067639, 0.00067609, 0.00067565, 
    0.00067511, 0.00067445, 0.00067361, 0.00067269, 0.00067149, 0.00067014, 
    0.00066856, 0.0006666, 0.00066446, 0.00066169, 0.00065865, 0.00065508, 
    0.00065079, 0.00064608, 0.00064012, 0.00063376, 0.0006266, 0.00061873, 
    0.00061035, 0.00060117, 0.00059183, 0.00058243, 0.00057345, 0.00056477, 
    0.00055684, 0.00054915, 0.00054229, 0.00053603, 0.00053035, 0.00052544, 
    0.0005207, 0.00051623, 0.00051195, 0.00050789, 0.00050418, 0.00050061, 
    0.00049752, 0.00049475, 0.00049243, 0.00049063, 0.00048905, 0.00048802, 
    0.00048721, 0.00048676, 0.00048659, 0.00048655, 0.00048655, 0.0004865, 
    0.00048638, 0.00048605, 0.00048561, 0.00048463, 0.00048339, 0.00048157, 
    0.00047919, 0.00047643, 0.00047281, 0.00046899, 0.00046482, 0.00046058, 
    0.00045627, 0.00045246, 0.00044884, 0.00044579, 0.00044307, 0.00044067, 
    0.00043878, 0.00043703, 0.00043552, 0.00043397, 0.00043236, 0.00043057, 
    0.00042874, 0.00042688, 0.00042494, 0.0004229, 0.00042078, 0.00041863, 
    0.00041639, 0.00041405, 0.00041153, 0.00040924, 0.00040704, 0.00040533, 
    0.0004036, 0.00040186, 0.00039992, 0.00039786, 0.00039561, 0.00039318, 
    0.00039034, 0.00038738, 0.00038433, 0.0003812, 0.00037799, 0.00037457, 
    0.00037099, 0.00036728, 0.00036334, 0.00035928, 0.00035497, 0.00035039, 
    0.00034554, 0.00034027, 0.00033478, 0.00032882, 0.00032271, 0.00031644, 
    0.0003103, 0.00030417, 0.00029831, 0.00029244, 0.00028657, 0.00028117, 
    0.00027592, 0.0002714, 0.00026715, 0.00026338, 0.00026018, 0.00025721, 
    0.00025467, 0.00025223, 0.00025001, 0.00024806, 0.00024624, 0.00024501, 
    0.00024389, 0.00024302, 0.00024245, 0.00024208, 0.00024184, 0.00024163, 
    0.00024152, 0.00024142, 0.00024135, 0.00024129, 0.00024123, 0.00024117, 
    0.0002411, 0.00024101, 0.0002409, 0.00024077, 0.0002406, 0.00024039, 
    0.00024016, 0.00023987, 0.00023957, 0.0002392, 0.00023883, 0.00023846, 
    0.00023811, 0.00023776, 0.00023739, 0.00023697, 0.0002365, 0.00023592, 
    0.00023528, 0.00023427, 0.00023309, 0.00023159, 0.0002297, 0.00022759, 
    0.00022486, 0.00022188, 0.00021835, 0.0002143, 0.00020987, 0.0002047, 
    0.00019921, 0.00019315, 0.00018684, 0.00018028, 0.000174, 0.00016771, 
    0.0001618, 0.00015609, 0.00015058, 0.00014558, 0.00014069, 0.00013645, 
    0.00013247, 0.00012882, 0.00012557, 0.00012243, 0.0001197, 0.00011704, 
    0.00011454, 0.00011208, 0.00010961, 0.00010711, 0.00010461, 0.00010217, 
    9.9813e-05, 9.7464e-05, 9.5672e-05, 9.4122e-05, 9.3106e-05, 9.2456e-05, 
    9.2005e-05, 9.1868e-05, 9.1786e-05, 9.1811e-05, 9.1838e-05, 9.1864e-05, 
    9.1774e-05, 9.1625e-05, 9.1318e-05, 9.0887e-05, 9.0356e-05, 8.976e-05, 
    8.9151e-05, 8.854e-05, 8.7933e-05, 8.7332e-05, 8.6748e-05, 8.6168e-05, 
    8.5609e-05, 8.5067e-05, 8.4546e-05, 8.4056e-05, 8.3578e-05, 8.3165e-05, 
    8.2796e-05, 8.2489e-05, 8.2334e-05, 8.2254e-05, 8.2502e-05, 8.2862e-05, 
    8.3406e-05, 8.4089e-05, 8.483e-05, 8.5637e-05, 8.6394e-05, 8.7058e-05, 
    8.7603e-05, 8.8083e-05, 8.839e-05, 8.8647e-05, 8.8793e-05, 8.8869e-05, 
    8.89e-05, 8.8833e-05, 8.8753e-05, 8.8657e-05, 8.857e-05, 8.8489e-05, 
    8.8384e-05, 8.8273e-05, 8.8146e-05, 8.8032e-05, 8.793e-05, 8.7849e-05, 
    8.7772e-05, 8.7699e-05, 8.7606e-05, 8.749e-05, 8.7289e-05, 8.7052e-05, 
    8.6715e-05, 8.6359e-05, 8.5979e-05, 8.5613e-05, 8.5255e-05, 8.4961e-05, 
    8.4718e-05, 8.4562e-05, 8.4534e-05, 8.4564e-05, 8.4755e-05, 8.4977e-05, 
    8.5259e-05, 8.5517e-05, 8.5762e-05, 8.5954e-05, 8.6133e-05, 8.6287e-05, 
    8.6417e-05, 8.653e-05, 8.6585e-05, 8.6622e-05, 8.6618e-05, 8.6572e-05, 
    8.6494e-05, 8.635e-05, 8.6198e-05, 8.6054e-05, 8.5909e-05, 8.5762e-05, 
    8.5583e-05, 8.5403e-05, 8.5253e-05, 8.5128e-05, 8.5032e-05, 8.4931e-05, 
    8.4825e-05, 8.4681e-05, 8.4524e-05, 8.4349e-05, 8.4124e-05, 8.3878e-05, 
    8.3596e-05, 8.3301e-05, 8.2984e-05, 8.2612e-05, 8.2214e-05, 8.1778e-05, 
    8.1345e-05, 8.0924e-05, 8.0576e-05, 8.0266e-05, 8.0095e-05, 7.9954e-05, 
    7.9875e-05, 7.9831e-05, 7.981e-05, 7.9809e-05, 7.9804e-05, 7.9783e-05, 
    7.9747e-05, 7.9698e-05, 7.9626e-05, 7.9545e-05, 7.9442e-05, 7.9339e-05, 
    7.9234e-05, 7.9118e-05, 7.8997e-05, 7.8872e-05, 7.8763e-05, 7.8672e-05, 
    7.86e-05, 7.8531e-05, 7.8442e-05, 7.8342e-05, 7.8227e-05, 7.8095e-05, 
    7.7954e-05, 7.7776e-05, 7.7583e-05, 7.7368e-05, 7.7104e-05, 7.6817e-05, 
    7.6465e-05, 7.6112e-05, 7.5758e-05, 7.5415e-05, 7.5079e-05, 7.4796e-05, 
    7.4529e-05, 7.4299e-05, 7.4098e-05, 7.3918e-05, 7.3795e-05, 7.369e-05, 
    7.363e-05, 7.3584e-05, 7.3551e-05, 7.3516e-05, 7.3479e-05, 7.3435e-05, 
    7.3386e-05, 7.3331e-05, 7.3254e-05, 7.3161e-05, 7.3013e-05, 7.284e-05, 
    7.2639e-05, 7.2415e-05, 7.2182e-05, 7.1927e-05, 7.1664e-05, 7.139e-05, 
    7.1119e-05, 7.085e-05, 7.0607e-05, 7.0388e-05, 7.0209e-05, 7.0071e-05, 
    6.9951e-05, 6.9874e-05, 6.9806e-05, 6.9753e-05, 6.9718e-05, 6.9692e-05, 
    6.9681e-05, 6.9672e-05, 6.9669e-05, 6.9666e-05, 6.9666e-05, 6.9663e-05, 
    6.9657e-05, 6.9644e-05, 6.9627e-05, 6.9607e-05, 6.9587e-05, 6.9568e-05, 
    6.9547e-05, 6.9525e-05, 6.9501e-05, 6.9477e-05, 6.9456e-05, 6.9446e-05, 
    6.9442e-05, 6.9445e-05, 6.9448e-05, 6.9452e-05, 6.9456e-05, 6.9461e-05, 
    6.9466e-05, 6.9471e-05, 6.9476e-05, 6.9484e-05, 6.9492e-05, 6.9504e-05, 
    6.9509e-05, 6.9511e-05, 6.9504e-05, 6.9498e-05, 6.9497e-05, 6.95e-05, 
    6.9507e-05, 6.9511e-05, 6.9513e-05, 6.9513e-05, 6.9512e-05, 6.9511e-05, 
    6.951e-05, 6.9515e-05, 6.9537e-05, 6.9572e-05, 6.9617e-05, 6.9663e-05, 
    6.9709e-05, 6.9753e-05, 6.9799e-05, 6.9848e-05, 6.9896e-05, 6.9941e-05, 
    6.9971e-05, 7.0001e-05, 7.0028e-05, 7.0051e-05, 7.0074e-05, 7.0111e-05, 
    7.0153e-05, 7.02e-05, 7.0258e-05, 7.032e-05, 7.0391e-05, 7.046e-05, 
    7.0525e-05, 7.0579e-05, 7.0627e-05, 7.0659e-05, 7.0683e-05, 7.0694e-05, 
    7.069e-05, 7.0679e-05, 7.0656e-05, 7.0623e-05, 7.0567e-05, 7.0493e-05, 
    7.0407e-05, 7.0313e-05, 7.0218e-05, 7.0127e-05, 7.0038e-05, 6.995e-05, 
    6.9848e-05, 6.9735e-05, 6.9594e-05, 6.9428e-05, 6.9238e-05, 6.8996e-05, 
    6.8731e-05, 6.8397e-05, 6.8019e-05, 6.7591e-05, 6.7099e-05, 6.6586e-05, 
    6.6053e-05, 6.5539e-05, 6.5051e-05, 6.4599e-05, 6.4163e-05, 6.38e-05, 
    6.3466e-05, 6.318e-05, 6.2935e-05, 6.2709e-05, 6.2538e-05, 6.2381e-05, 
    6.2251e-05, 6.2132e-05, 6.2019e-05, 6.192e-05, 6.183e-05, 6.176e-05, 
    6.1708e-05, 6.1667e-05, 6.1644e-05, 6.1623e-05, 6.1609e-05, 6.1594e-05, 
    6.1578e-05, 6.1563e-05, 6.1549e-05, 6.1542e-05, 6.1539e-05, 6.154e-05, 
    6.154e-05, 6.1539e-05, 6.153e-05, 6.1511e-05, 6.148e-05, 6.1428e-05, 
    6.1367e-05, 6.1284e-05, 6.1197e-05, 6.1103e-05, 6.1003e-05, 6.0903e-05, 
    6.0816e-05, 6.0735e-05, 6.0662e-05, 6.0595e-05, 6.0531e-05, 6.0472e-05, 
    6.0415e-05, 6.036e-05, 6.0302e-05, 6.0242e-05, 6.0166e-05, 6.0089e-05, 
    6.0009e-05, 5.9926e-05, 5.9842e-05, 5.9752e-05, 5.9661e-05, 5.9567e-05, 
    5.9473e-05, 5.9378e-05, 5.9289e-05, 5.9205e-05, 5.914e-05, 5.9086e-05, 
    5.9044e-05, 5.9014e-05, 5.8989e-05, 5.8975e-05, 5.8964e-05, 5.8957e-05, 
    5.8954e-05, 5.8951e-05, 5.8951e-05, 5.8948e-05, 5.8944e-05, 5.8938e-05, 
    5.8932e-05, 5.8919e-05, 5.8902e-05, 5.8877e-05, 5.8841e-05, 5.8799e-05, 
    5.8737e-05, 5.8667e-05, 5.8583e-05, 5.8487e-05, 5.8386e-05, 5.827e-05, 
    5.8156e-05, 5.8047e-05, 5.7958e-05, 5.7881e-05, 5.7846e-05, 5.7822e-05, 
    5.7818e-05, 5.7815e-05, 5.7813e-05, 5.7792e-05, 5.7765e-05, 5.772e-05, 
    5.7669e-05, 5.7613e-05, 5.7553e-05, 5.7494e-05, 5.7447e-05, 5.7416e-05, 
    5.7401e-05, 5.7405e-05, 5.7415e-05, 5.7436e-05, 5.7458e-05, 5.748e-05, 
    5.7493e-05, 5.7503e-05, 5.7504e-05, 5.7506e-05, 5.7511e-05, 5.7522e-05, 
    5.7535e-05, 5.7516e-05, 5.7462e-05, 5.734e-05, 5.7114e-05, 5.6831e-05, 
    5.6318e-05, 5.5703e-05, 5.4859e-05, 5.3839e-05, 5.2692e-05, 5.1357e-05, 
    4.9968e-05, 4.8521e-05, 4.7193e-05, 4.5957e-05, 4.4988e-05, 4.4096e-05, 
    4.3422e-05, 4.2866e-05, 4.2426e-05, 4.2136e-05, 4.1894e-05, 4.1762e-05, 
    4.166e-05, 4.159e-05, 4.1539e-05, 4.1492e-05, 4.1439e-05, 4.1379e-05, 
    4.1306e-05, 4.118e-05, 4.1029e-05, 4.0787e-05, 4.0505e-05, 4.0158e-05, 
    3.9831e-05, 3.9515e-05, 3.9383e-05, 3.9307e-05, 3.9344e-05, 3.9457e-05, 
    3.9611e-05, 3.9786e-05, 3.9939e-05, 4.0037e-05, 4.0038e-05, 3.9978e-05, 
    3.972e-05, 3.9391e-05, 3.8885e-05, 3.8295e-05, 3.7634e-05, 3.701e-05, 
    3.6399e-05, 3.5855e-05, 3.5345e-05, 3.4869e-05, 3.4452e-05, 3.4058e-05, 
    3.3741e-05, 3.3469e-05, 3.3247e-05, 3.3074e-05, 3.292e-05, 3.2821e-05, 
    3.2746e-05, 3.2703e-05, 3.2682e-05, 3.2669e-05, 3.2665e-05, 3.2661e-05, 
    3.2659e-05, 3.2654e-05, 3.2647e-05, 3.2642e-05, 3.2642e-05, 3.2649e-05, 
    3.2662e-05, 3.2678e-05, 3.2695e-05, 3.2711e-05, 3.2724e-05, 3.274e-05, 
    3.2756e-05, 3.2778e-05, 3.28e-05, 3.282e-05, 3.2842e-05, 3.2866e-05, 
    3.2886e-05, 3.2905e-05, 3.2922e-05, 3.2937e-05, 3.295e-05, 3.2961e-05, 
    3.297e-05, 3.2973e-05, 3.2975e-05, 3.2976e-05, 3.2977e-05, 3.2977e-05, 
    3.2975e-05, 3.2973e-05, 3.2971e-05, 3.297e-05, 3.297e-05, 3.2972e-05, 
    3.2973e-05, 3.2975e-05, 3.2975e-05, 3.2974e-05, 3.2976e-05, 3.2977e-05, 
    3.2976e-05, 3.2962e-05, 3.2942e-05, 3.2908e-05, 3.2874e-05, 3.284e-05, 
    3.2818e-05, 3.2803e-05, 3.2805e-05, 3.2809e-05, 3.2819e-05, 3.283e-05, 
    3.2842e-05, 3.2866e-05, 3.2891e-05, 3.2919e-05, 3.2944e-05, 3.2965e-05, 
    3.2984e-05, 3.3005e-05, 3.3035e-05, 3.3059e-05, 3.3079e-05, 3.3093e-05, 
    3.3104e-05, 3.3115e-05, 3.3124e-05, 3.313e-05, 3.3135e-05, 3.3138e-05, 
    3.3146e-05, 3.3156e-05, 3.3169e-05, 3.3184e-05, 3.3202e-05, 3.3226e-05, 
    3.3251e-05, 3.3279e-05, 3.3306e-05, 3.3331e-05, 3.3356e-05, 3.3381e-05, 
    3.3407e-05, 3.3433e-05, 3.3458e-05, 3.3486e-05, 3.3513e-05, 3.3535e-05, 
    3.3553e-05, 3.3565e-05, 3.3564e-05, 3.356e-05, 3.3551e-05, 3.3544e-05, 
    3.3539e-05, 3.3537e-05, 3.3535e-05, 3.3529e-05, 3.3521e-05, 3.3512e-05, 
    3.3502e-05, 3.3492e-05, 3.3487e-05, 3.3484e-05, 3.3481e-05, 3.3483e-05, 
    3.3487e-05, 3.3496e-05, 3.3505e-05, 3.3514e-05, 3.3523e-05, 3.3533e-05, 
    3.3548e-05, 3.3566e-05, 3.359e-05, 3.3617e-05, 3.3647e-05, 3.369e-05, 
    3.3732e-05, 3.3767e-05, 3.3785e-05, 3.3792e-05, 3.38e-05, 3.381e-05, 
    3.3823e-05, 3.3823e-05, 3.3814e-05, 3.3786e-05, 3.3752e-05, 3.3707e-05, 
    3.3648e-05, 3.3578e-05, 3.3486e-05, 3.3389e-05, 3.3286e-05, 3.3171e-05, 
    3.3043e-05, 3.2895e-05, 3.2738e-05, 3.2562e-05, 3.2377e-05, 3.2183e-05, 
    3.1978e-05, 3.177e-05, 3.1566e-05, 3.1377e-05, 3.1213e-05, 3.1052e-05, 
    3.0892e-05, 3.0741e-05, 3.0588e-05, 3.0433e-05, 3.029e-05, 3.0154e-05, 
    3.0007e-05, 2.9854e-05, 2.9686e-05, 2.9524e-05, 2.9366e-05, 2.9234e-05, 
    2.9105e-05, 2.8982e-05, 2.8874e-05, 2.8778e-05, 2.8726e-05, 2.8685e-05, 
    2.8666e-05, 2.8662e-05, 2.8673e-05, 2.871e-05, 2.8757e-05, 2.8819e-05, 
    2.8878e-05, 2.8931e-05, 2.8984e-05, 2.9037e-05, 2.9083e-05, 2.9114e-05, 
    2.9125e-05, 2.9102e-05, 2.9065e-05, 2.9007e-05, 2.8944e-05, 2.887e-05, 
    2.8792e-05, 2.871e-05, 2.8619e-05, 2.8529e-05, 2.844e-05, 2.8364e-05, 
    2.8296e-05, 2.8244e-05, 2.8194e-05, 2.8149e-05, 2.8115e-05, 2.8088e-05, 
    2.8076e-05, 2.8067e-05, 2.8061e-05, 2.8061e-05, 2.8066e-05, 2.8074e-05, 
    2.8083e-05, 2.8097e-05, 2.811e-05, 2.8124e-05, 2.8144e-05, 2.8165e-05, 
    2.8185e-05, 2.8203e-05, 2.8218e-05, 2.8234e-05, 2.8251e-05, 2.8273e-05, 
    2.8294e-05, 2.8316e-05, 2.8342e-05, 2.837e-05, 2.8401e-05, 2.843e-05, 
    2.8456e-05, 2.8479e-05, 2.8499e-05, 2.8495e-05, 2.8487e-05, 2.8473e-05, 
    2.8451e-05, 2.8425e-05, 2.8404e-05, 2.8378e-05, 2.834e-05, 2.8308e-05, 
    2.8279e-05, 2.8257e-05, 2.8237e-05, 2.822e-05, 2.8203e-05, 2.8186e-05, 
    2.8168e-05, 2.815e-05, 2.8131e-05, 2.8115e-05, 2.8103e-05, 2.8097e-05, 
    2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8092e-05, 2.8093e-05, 
    2.81e-05, 2.8111e-05, 2.8128e-05, 2.8147e-05, 2.8168e-05, 2.8215e-05, 
    2.8271e-05, 2.834e-05, 2.8425e-05, 2.8516e-05, 2.8617e-05, 2.8712e-05, 
    2.88e-05, 2.887e-05, 2.8931e-05, 2.8979e-05, 2.9025e-05, 2.9069e-05, 
    2.9106e-05, 2.9137e-05, 2.9163e-05, 2.9186e-05, 2.9206e-05, 2.9226e-05, 
    2.9245e-05, 2.9265e-05, 2.9286e-05, 2.9308e-05, 2.9328e-05, 2.9348e-05, 
    2.9366e-05, 2.9382e-05, 2.9396e-05, 2.9412e-05, 2.9431e-05, 2.9455e-05, 
    2.948e-05, 2.9504e-05, 2.9527e-05, 2.9548e-05, 2.9566e-05, 2.9583e-05, 
    2.9603e-05, 2.9622e-05, 2.9637e-05, 2.9653e-05, 2.967e-05, 2.9678e-05, 
    2.9683e-05, 2.9685e-05, 2.9688e-05, 2.969e-05, 2.9706e-05, 2.9722e-05, 
    2.9736e-05, 2.9753e-05, 2.9771e-05, 2.9795e-05, 2.982e-05, 2.9848e-05, 
    2.9878e-05, 2.991e-05, 2.9947e-05, 2.9987e-05, 3.0027e-05, 3.0064e-05, 
    3.0099e-05, 3.0126e-05, 3.0152e-05, 3.0173e-05, 3.0193e-05, 3.0212e-05, 
    3.0223e-05, 3.023e-05, 3.0226e-05, 3.0214e-05, 3.0193e-05, 3.0153e-05, 
    3.0105e-05, 3.0043e-05, 2.997e-05, 2.9881e-05, 2.9778e-05, 2.9669e-05, 
    2.954e-05, 2.9406e-05, 2.9264e-05, 2.9103e-05, 2.8933e-05, 2.8747e-05, 
    2.8548e-05, 2.8321e-05, 2.8073e-05, 2.781e-05, 2.7528e-05, 2.7246e-05, 
    2.6973e-05, 2.6698e-05, 2.6424e-05, 2.6148e-05, 2.5875e-05, 2.5614e-05, 
    2.5371e-05, 2.5144e-05, 2.4953e-05, 2.4774e-05, 2.4626e-05, 2.4484e-05, 
    2.435e-05, 2.4189e-05, 2.4022e-05, 2.3855e-05, 2.3698e-05, 2.3555e-05, 
    2.3427e-05, 2.3305e-05, 2.3202e-05, 2.3101e-05, 2.3001e-05, 2.2912e-05, 
    2.2828e-05, 2.2745e-05, 2.2667e-05, 2.2602e-05, 2.255e-05, 2.2505e-05, 
    2.2452e-05, 2.2401e-05, 2.2351e-05, 2.2313e-05, 2.2282e-05, 2.2258e-05, 
    2.2234e-05, 2.2208e-05, 2.2186e-05, 2.2166e-05, 2.2147e-05, 2.213e-05, 
    2.212e-05, 2.2115e-05, 2.2115e-05, 2.2113e-05, 2.211e-05, 2.2105e-05, 
    2.2104e-05, 2.2107e-05, 2.211e-05, 2.2113e-05, 2.2112e-05, 2.2111e-05, 
    2.2108e-05, 2.2108e-05, 2.2109e-05, 2.2109e-05, 2.2112e-05, 2.2117e-05, 
    2.2122e-05, 2.2125e-05, 2.2125e-05, 2.2125e-05, 2.2126e-05, 2.2125e-05, 
    2.2125e-05, 2.2125e-05, 2.2126e-05, 2.213e-05, 2.2139e-05, 2.2152e-05, 
    2.2176e-05, 2.2199e-05, 2.2217e-05, 2.2228e-05, 2.2234e-05, 2.2243e-05, 
    2.2253e-05, 2.2268e-05, 2.2283e-05, 2.2299e-05, 2.2313e-05, 2.2327e-05, 
    2.2339e-05, 2.2352e-05, 2.2366e-05, 2.2376e-05, 2.2382e-05, 2.2372e-05, 
    2.2355e-05, 2.2329e-05, 2.2298e-05, 2.2265e-05, 2.2227e-05, 2.2184e-05, 
    2.2134e-05, 2.2094e-05, 2.2059e-05, 2.2031e-05, 2.2002e-05, 2.1972e-05, 
    2.1947e-05, 2.1926e-05, 2.1913e-05, 2.1901e-05, 2.1887e-05, 2.187e-05, 
    2.185e-05, 2.1823e-05, 2.1795e-05, 2.1761e-05, 2.1728e-05, 2.1694e-05, 
    2.1667e-05, 2.1641e-05, 2.1616e-05, 2.1586e-05, 2.155e-05, 2.1509e-05, 
    2.1466e-05, 2.1427e-05, 2.1389e-05, 2.1355e-05, 2.1324e-05, 2.1295e-05, 
    2.1274e-05, 2.1257e-05, 2.1246e-05, 2.124e-05, 2.1236e-05, 2.1238e-05, 
    2.1243e-05, 2.1251e-05, 2.1262e-05, 2.1274e-05, 2.129e-05, 2.1305e-05, 
    2.1321e-05, 2.1339e-05, 2.1358e-05, 2.1377e-05, 2.1392e-05, 2.1397e-05, 
    2.1399e-05, 2.1398e-05, 2.1393e-05, 2.1385e-05, 2.1367e-05, 2.1343e-05, 
    2.1313e-05, 2.1272e-05, 2.1226e-05, 2.1162e-05, 2.1098e-05, 2.1031e-05, 
    2.098e-05, 2.0931e-05, 2.0875e-05, 2.0814e-05, 2.0747e-05, 2.0687e-05, 
    2.063e-05, 2.0594e-05, 2.0562e-05, 2.0535e-05, 2.0519e-05, 2.0507e-05, 
    2.0508e-05, 2.0505e-05, 2.0498e-05, 2.0484e-05, 2.0466e-05, 2.0439e-05, 
    2.0413e-05, 2.0386e-05, 2.035e-05, 2.0308e-05, 2.0288e-05, 2.0272e-05, 
    2.0263e-05, 2.0254e-05, 2.0245e-05, 2.0236e-05, 2.0228e-05, 2.0226e-05, 
    2.0235e-05, 2.0251e-05, 2.0297e-05, 2.0352e-05, 2.0429e-05, 2.0531e-05, 
    2.0656e-05, 2.0826e-05, 2.1016e-05, 2.1268e-05, 2.1561e-05, 2.1897e-05, 
    2.2239e-05, 2.2577e-05, 2.2895e-05, 2.3225e-05, 2.3571e-05, 2.3945e-05, 
    2.4323e-05, 2.4676e-05, 2.5003e-05, 2.5292e-05, 2.5555e-05, 2.5803e-05, 
    2.6005e-05, 2.6193e-05, 2.6352e-05, 2.6499e-05, 2.664e-05, 2.677e-05, 
    2.6892e-05, 2.6995e-05, 2.7091e-05, 2.7182e-05, 2.727e-05, 2.7354e-05, 
    2.7428e-05, 2.7495e-05, 2.7557e-05, 2.7599e-05, 2.7634e-05, 2.7653e-05, 
    2.7671e-05, 2.7688e-05, 2.7698e-05, 2.7707e-05, 2.7711e-05, 2.7718e-05, 
    2.7728e-05, 2.7738e-05, 2.7749e-05, 2.7765e-05, 2.7783e-05, 2.7802e-05, 
    2.7824e-05, 2.7846e-05, 2.786e-05, 2.7874e-05, 2.7887e-05, 2.7897e-05, 
    2.7905e-05, 2.7907e-05, 2.7905e-05, 2.7894e-05, 2.7882e-05, 2.7869e-05, 
    2.7847e-05, 2.782e-05, 2.7785e-05, 2.7749e-05, 2.7714e-05, 2.7682e-05, 
    2.7655e-05, 2.764e-05, 2.7631e-05, 2.7627e-05, 2.7628e-05, 2.763e-05, 
    2.7639e-05, 2.7654e-05, 2.7676e-05, 2.7712e-05, 2.7756e-05, 2.7818e-05, 
    2.789e-05, 2.7972e-05, 2.8074e-05, 2.8183e-05, 2.8306e-05, 2.8425e-05, 
    2.854e-05, 2.8642e-05, 2.8738e-05, 2.881e-05, 2.8874e-05, 2.8924e-05, 
    2.8962e-05, 2.8994e-05, 2.9014e-05, 2.9028e-05, 2.903e-05, 2.9021e-05, 
    2.9005e-05, 2.8987e-05, 2.8961e-05, 2.8918e-05, 2.8865e-05, 2.8805e-05, 
    2.8735e-05, 2.8666e-05, 2.8606e-05, 2.8567e-05, 2.8544e-05, 2.8571e-05, 
    2.8614e-05, 2.8693e-05, 2.879e-05, 2.8904e-05, 2.9042e-05, 2.9187e-05, 
    2.9344e-05, 2.9498e-05, 2.9651e-05, 2.9789e-05, 2.9922e-05, 3.0038e-05, 
    3.0143e-05, 3.0235e-05, 3.031e-05, 3.0378e-05, 3.0427e-05, 3.0469e-05, 
    3.0498e-05, 3.0512e-05, 3.0519e-05, 3.0509e-05, 3.0497e-05, 3.0479e-05, 
    3.0455e-05, 3.0428e-05, 3.0396e-05, 3.0361e-05, 3.0316e-05, 3.0274e-05, 
    3.0233e-05, 3.0186e-05, 3.0143e-05, 3.0109e-05, 3.0081e-05, 3.0056e-05, 
    3.0046e-05, 3.0039e-05, 3.0039e-05, 3.004e-05, 3.0043e-05, 3.0045e-05, 
    3.0046e-05, 3.0043e-05, 3.0037e-05, 3.0025e-05, 3.0004e-05, 2.9979e-05, 
    2.9948e-05, 2.9916e-05, 2.988e-05, 2.9847e-05, 2.9814e-05, 2.9788e-05, 
    2.9763e-05, 2.9738e-05, 2.9716e-05, 2.9695e-05, 2.9685e-05, 2.9677e-05, 
    2.9676e-05, 2.968e-05, 2.9688e-05, 2.9706e-05, 2.9726e-05, 2.9751e-05, 
    2.9782e-05, 2.9817e-05, 2.9856e-05, 2.9894e-05, 2.9928e-05, 2.9957e-05, 
    2.9982e-05, 2.9998e-05, 3.0013e-05, 3.0028e-05, 3.004e-05, 3.0048e-05, 
    3.0054e-05, 3.0058e-05, 3.0061e-05, 3.0062e-05, 3.0062e-05, 3.006e-05, 
    3.0057e-05, 3.0052e-05, 3.0045e-05, 3.0036e-05, 3.0022e-05, 3.0007e-05, 
    2.9987e-05, 2.9965e-05, 2.9938e-05, 2.9909e-05, 2.9879e-05, 2.9856e-05, 
    2.9837e-05, 2.9824e-05, 2.9814e-05, 2.9804e-05, 2.9796e-05, 2.9789e-05, 
    2.978e-05, 2.9779e-05, 2.9782e-05, 2.9801e-05, 2.9823e-05, 2.9854e-05, 
    2.9881e-05, 2.9905e-05, 2.9912e-05, 2.9916e-05, 2.992e-05, 2.9923e-05, 
    2.9925e-05, 2.9924e-05, 2.9921e-05, 2.9918e-05, 2.9918e-05, 2.9922e-05, 
    2.9928e-05, 2.9934e-05, 2.9938e-05, 2.9938e-05, 2.9935e-05, 2.993e-05, 
    2.9924e-05, 2.9916e-05, 2.9909e-05, 2.9904e-05, 2.9899e-05, 2.9894e-05, 
    2.9881e-05, 2.9872e-05, 2.9869e-05, 2.9872e-05, 2.9878e-05, 2.9892e-05, 
    2.9904e-05, 2.9913e-05, 2.9918e-05, 2.9921e-05, 2.9926e-05, 2.9932e-05, 
    2.9943e-05, 2.9958e-05, 2.9976e-05, 2.9986e-05, 2.9995e-05, 2.9997e-05, 
    2.9997e-05, 2.9993e-05, 2.9981e-05, 2.9968e-05, 2.9948e-05, 2.9932e-05, 
    2.992e-05, 2.9922e-05, 2.9929e-05, 2.9941e-05, 2.995e-05, 2.9956e-05, 
    2.9957e-05, 2.9957e-05, 2.996e-05, 2.9964e-05, 2.9969e-05, 2.9973e-05, 
    2.9977e-05, 2.9984e-05, 2.9989e-05, 2.9988e-05, 2.9991e-05, 2.9996e-05, 
    3.0011e-05, 3.0031e-05, 3.0063e-05, 3.0092e-05, 3.0121e-05, 3.0134e-05, 
    3.0144e-05, 3.0146e-05, 3.0146e-05, 3.0145e-05, 3.0143e-05, 3.0142e-05, 
    3.014e-05, 3.0141e-05, 3.0143e-05, 3.015e-05, 3.016e-05, 3.0175e-05, 
    3.0191e-05, 3.0208e-05, 3.0223e-05, 3.0236e-05, 3.0244e-05, 3.0251e-05, 
    3.0255e-05, 3.0257e-05, 3.0258e-05, 3.0256e-05, 3.0253e-05, 3.0249e-05, 
    3.0244e-05, 3.024e-05, 3.0244e-05, 3.0251e-05, 3.0267e-05, 3.0294e-05, 
    3.0325e-05, 3.0345e-05, 3.0365e-05, 3.0389e-05, 3.0419e-05, 3.0455e-05, 
    3.0504e-05, 3.0557e-05, 3.0615e-05, 3.0684e-05, 3.0761e-05, 3.0862e-05, 
    3.0971e-05, 3.1098e-05, 3.1242e-05, 3.14e-05, 3.1585e-05, 3.1777e-05, 
    3.1979e-05, 3.2181e-05, 3.2385e-05, 3.2562e-05, 3.2729e-05, 3.2876e-05, 
    3.3014e-05, 3.3138e-05, 3.3259e-05, 3.3378e-05, 3.3497e-05, 3.3616e-05, 
    3.3734e-05, 3.3837e-05, 3.3933e-05, 3.3999e-05, 3.4055e-05, 3.4092e-05, 
    3.4117e-05, 3.4136e-05, 3.4156e-05, 3.4179e-05, 3.4208e-05, 3.4225e-05, 
    3.4236e-05, 3.4237e-05, 3.4238e-05, 3.4239e-05, 3.4242e-05, 3.4247e-05, 
    3.4253e-05, 3.4258e-05, 3.4262e-05, 3.4265e-05, 3.4266e-05, 3.4265e-05, 
    3.4263e-05, 3.426e-05, 3.4255e-05, 3.4248e-05, 3.4235e-05, 3.4219e-05, 
    3.4188e-05, 3.4151e-05, 3.4106e-05, 3.404e-05, 3.3963e-05, 3.3853e-05, 
    3.3724e-05, 3.3562e-05, 3.3357e-05, 3.3132e-05, 3.2897e-05, 3.266e-05, 
    3.2425e-05, 3.2164e-05, 3.1889e-05, 3.1571e-05, 3.125e-05, 3.0926e-05, 
    3.0619e-05, 3.0322e-05, 3.0058e-05, 2.9802e-05, 2.9567e-05, 2.935e-05, 
    2.9146e-05, 2.8969e-05, 2.8801e-05, 2.8658e-05, 2.8529e-05, 2.8414e-05, 
    2.8318e-05, 2.8227e-05, 2.8142e-05, 2.8063e-05, 2.7989e-05, 2.7917e-05, 
    2.7847e-05, 2.7783e-05, 2.7725e-05, 2.7672e-05, 2.762e-05, 2.7569e-05, 
    2.7521e-05, 2.7471e-05, 2.7417e-05, 2.736e-05, 2.7302e-05, 2.7245e-05, 
    2.7189e-05, 2.7135e-05, 2.7078e-05, 2.7021e-05, 2.6967e-05, 2.6914e-05, 
    2.6866e-05, 2.6824e-05, 2.6785e-05, 2.6757e-05, 2.6732e-05, 2.6713e-05, 
    2.6697e-05, 2.6685e-05, 2.6675e-05, 2.6665e-05, 2.6658e-05, 2.6652e-05, 
    2.6647e-05, 2.6644e-05, 2.6641e-05, 2.664e-05, 2.6642e-05, 2.6649e-05, 
    2.6658e-05, 2.6669e-05, 2.6677e-05, 2.6684e-05, 2.6687e-05, 2.6686e-05, 
    2.6682e-05, 2.6656e-05, 2.6618e-05, 2.656e-05, 2.6479e-05, 2.6387e-05, 
    2.6269e-05, 2.6145e-05, 2.6011e-05, 2.5883e-05, 2.5759e-05, 2.5654e-05, 
    2.5559e-05, 2.5486e-05, 2.5433e-05, 2.5394e-05, 2.5385e-05, 2.5381e-05, 
    2.5387e-05, 2.5401e-05, 2.5421e-05, 2.5453e-05, 2.5488e-05, 2.553e-05, 
    2.5569e-05, 2.5606e-05, 2.5635e-05, 2.5661e-05, 2.5674e-05, 2.5681e-05, 
    2.5681e-05, 2.5658e-05, 2.5625e-05, 2.5558e-05, 2.5473e-05, 2.5366e-05, 
    2.5239e-05, 2.5105e-05, 2.4962e-05, 2.4813e-05, 2.4654e-05, 2.4487e-05, 
    2.4315e-05, 2.4147e-05, 2.3982e-05, 2.3827e-05, 2.3691e-05, 2.3566e-05, 
    2.348e-05, 2.3402e-05, 2.3342e-05, 2.3297e-05, 2.3262e-05, 2.324e-05, 
    2.3222e-05, 2.3211e-05, 2.3209e-05, 2.3212e-05, 2.3219e-05, 2.3227e-05, 
    2.3232e-05, 2.3236e-05, 2.3237e-05, 2.3236e-05, 2.3233e-05, 2.3227e-05, 
    2.3217e-05, 2.3202e-05, 2.3178e-05, 2.3148e-05, 2.31e-05, 2.3046e-05, 
    2.2981e-05, 2.2914e-05, 2.2845e-05, 2.2779e-05, 2.2717e-05, 2.2662e-05, 
    2.2623e-05, 2.259e-05, 2.2585e-05, 2.2587e-05, 2.2603e-05, 2.2624e-05, 
    2.2648e-05, 2.2664e-05, 2.2676e-05, 2.268e-05, 2.2682e-05, 2.2682e-05, 
    2.2682e-05, 2.2683e-05, 2.2688e-05, 2.2701e-05, 2.2719e-05, 2.2744e-05, 
    2.2767e-05, 2.2781e-05, 2.2782e-05, 2.2773e-05, 2.274e-05, 2.27e-05, 
    2.2648e-05, 2.26e-05, 2.2555e-05, 2.2517e-05, 2.2482e-05, 2.2461e-05, 
    2.2439e-05, 2.2416e-05, 2.2401e-05, 2.2389e-05, 2.2383e-05, 2.238e-05, 
    2.238e-05, 2.2384e-05, 2.239e-05, 2.2401e-05, 2.2413e-05, 2.2427e-05, 
    2.2439e-05, 2.245e-05, 2.2455e-05, 2.2457e-05, 2.2454e-05, 2.245e-05, 
    2.2445e-05, 2.2443e-05, 2.2443e-05, 2.2446e-05, 2.2454e-05, 2.2464e-05, 
    2.248e-05, 2.2496e-05, 2.2516e-05, 2.2536e-05, 2.2555e-05, 2.2568e-05, 
    2.2577e-05, 2.2563e-05, 2.2543e-05, 2.2517e-05, 2.2495e-05, 2.2474e-05, 
    2.2464e-05, 2.2458e-05, 2.2455e-05, 2.2455e-05, 2.2456e-05, 2.2459e-05, 
    2.2461e-05, 2.2462e-05, 2.2459e-05, 2.2453e-05, 2.2448e-05, 2.2443e-05, 
    2.2438e-05, 2.2435e-05, 2.2432e-05, 2.2429e-05, 2.2424e-05, 2.2416e-05, 
    2.2402e-05, 2.2383e-05, 2.2359e-05, 2.2335e-05, 2.2316e-05, 2.2294e-05, 
    2.2269e-05, 2.2238e-05, 2.2205e-05, 2.2164e-05, 2.213e-05, 2.2102e-05, 
    2.2085e-05, 2.207e-05, 2.206e-05, 2.2047e-05, 2.2031e-05, 2.2009e-05, 
    2.1986e-05, 2.1973e-05, 2.1963e-05, 2.1959e-05, 2.1958e-05, 2.1958e-05, 
    2.1958e-05, 2.1959e-05, 2.196e-05, 2.1957e-05, 2.1952e-05, 2.1937e-05, 
    2.1923e-05, 2.1914e-05, 2.1907e-05, 2.1901e-05, 2.1909e-05, 2.192e-05, 
    2.1935e-05, 2.1944e-05, 2.1951e-05, 2.1951e-05, 2.1948e-05, 2.1943e-05, 
    2.1945e-05, 2.1953e-05, 2.1962e-05, 2.197e-05, 2.1974e-05, 2.1976e-05, 
    2.1975e-05, 2.1992e-05, 2.2018e-05, 2.2073e-05, 2.2142e-05, 2.2225e-05, 
    2.2329e-05, 2.2441e-05, 2.2578e-05, 2.2726e-05, 2.2888e-05, 2.3047e-05, 
    2.3203e-05, 2.3333e-05, 2.3459e-05, 2.3579e-05, 2.37e-05, 2.3819e-05, 
    2.3927e-05, 2.4028e-05, 2.4114e-05, 2.4197e-05, 2.4278e-05, 2.4367e-05, 
    2.4463e-05, 2.4573e-05, 2.4695e-05, 2.4825e-05, 2.496e-05, 2.5091e-05, 
    2.5212e-05, 2.5324e-05, 2.543e-05, 2.5523e-05, 2.562e-05, 2.5737e-05, 
    2.5849e-05, 2.5956e-05, 2.6041e-05, 2.6118e-05, 2.6175e-05, 2.6222e-05, 
    2.6258e-05, 2.6261e-05, 2.6247e-05, 2.6175e-05, 2.6083e-05, 2.5962e-05, 
    2.58e-05, 2.5619e-05, 2.5387e-05, 2.5141e-05, 2.4874e-05, 2.4595e-05, 
    2.4311e-05, 2.4063e-05, 2.3822e-05, 2.3595e-05, 2.3387e-05, 2.3189e-05, 
    2.3004e-05, 2.282e-05, 2.2636e-05, 2.2455e-05, 2.2277e-05, 2.2126e-05, 
    2.1988e-05, 2.1886e-05, 2.1807e-05, 2.1746e-05, 2.1698e-05, 2.1651e-05, 
    2.1599e-05, 2.1542e-05, 2.148e-05, 2.1449e-05, 2.1428e-05, 2.1432e-05, 
    2.1445e-05, 2.1466e-05, 2.1497e-05, 2.153e-05, 2.1565e-05, 2.16e-05, 
    2.1634e-05, 2.1678e-05, 2.1727e-05, 2.179e-05, 2.185e-05, 2.1902e-05, 
    2.1933e-05, 2.1953e-05, 2.1959e-05, 2.1965e-05, 2.1969e-05, 2.1978e-05, 
    2.1988e-05, 2.2003e-05, 2.2017e-05, 2.2027e-05, 2.2032e-05, 2.2035e-05, 
    2.2037e-05, 2.2039e-05, 2.2042e-05, 2.2046e-05, 2.2052e-05, 2.2058e-05, 
    2.2062e-05, 2.2065e-05, 2.2066e-05, 2.2067e-05, 2.2067e-05, 2.2067e-05, 
    2.207e-05, 2.2074e-05, 2.2079e-05, 2.2084e-05, 2.2088e-05, 2.209e-05, 
    2.209e-05, 2.2089e-05, 2.2086e-05, 2.2083e-05, 2.2081e-05, 2.2085e-05, 
    2.2096e-05, 2.2113e-05, 2.2133e-05, 2.2155e-05, 2.2179e-05, 2.2204e-05, 
    2.2232e-05, 2.2262e-05, 2.2299e-05, 2.2336e-05, 2.2369e-05, 2.2393e-05, 
    2.241e-05, 2.2417e-05, 2.2424e-05, 2.2427e-05, 2.2428e-05, 2.2428e-05, 
    2.2428e-05, 2.2427e-05, 2.2427e-05, 2.2426e-05, 2.2426e-05, 2.2427e-05, 
    2.2427e-05, 2.2427e-05, 2.2429e-05, 2.2433e-05, 2.244e-05, 2.2447e-05, 
    2.2454e-05, 2.246e-05, 2.2464e-05, 2.2467e-05, 2.247e-05, 2.2472e-05, 
    2.2474e-05, 2.2477e-05, 2.2475e-05, 2.247e-05, 2.2462e-05, 2.2456e-05, 
    2.2451e-05, 2.2443e-05, 2.2435e-05, 2.2419e-05, 2.2402e-05, 2.2387e-05, 
    2.238e-05, 2.238e-05, 2.2399e-05, 2.2423e-05, 2.2457e-05, 2.2503e-05, 
    2.2559e-05, 2.263e-05, 2.2705e-05, 2.2791e-05, 2.2875e-05, 2.2957e-05, 
    2.3022e-05, 2.3081e-05, 2.3122e-05, 2.3156e-05, 2.3183e-05, 2.3208e-05, 
    2.3232e-05, 2.3253e-05, 2.3272e-05, 2.329e-05, 2.3318e-05, 2.335e-05, 
    2.3391e-05, 2.3434e-05, 2.3478e-05, 2.3504e-05, 2.3524e-05, 2.3524e-05, 
    2.3522e-05, 2.3515e-05, 2.3503e-05, 2.3488e-05, 2.3456e-05, 2.3419e-05, 
    2.3372e-05, 2.3329e-05, 2.3288e-05, 2.3267e-05, 2.3253e-05, 2.3254e-05, 
    2.3258e-05, 2.3264e-05, 2.3259e-05, 2.325e-05, 2.3226e-05, 2.3203e-05, 
    2.318e-05, 2.3162e-05, 2.3147e-05, 2.3141e-05, 2.3138e-05, 2.3138e-05, 
    2.3136e-05, 2.3133e-05, 2.3131e-05, 2.3131e-05, 2.3135e-05, 2.3147e-05, 
    2.3161e-05, 2.3174e-05, 2.3185e-05, 2.3193e-05, 2.3198e-05, 2.3202e-05, 
    2.3206e-05, 2.321e-05, 2.3218e-05, 2.3227e-05, 2.3238e-05, 2.3246e-05, 
    2.3252e-05, 2.3254e-05, 2.3252e-05, 2.3246e-05, 2.323e-05, 2.321e-05, 
    2.3183e-05, 2.315e-05, 2.3114e-05, 2.3085e-05, 2.3061e-05, 2.3051e-05, 
    2.3047e-05, 2.3049e-05, 2.3053e-05, 2.3057e-05, 2.3062e-05, 2.3062e-05, 
    2.306e-05, 2.3044e-05, 2.3024e-05, 2.2989e-05, 2.2956e-05, 2.2924e-05, 
    2.2904e-05, 2.289e-05, 2.2896e-05, 2.2905e-05, 2.2917e-05, 2.2927e-05, 
    2.2937e-05, 2.2945e-05, 2.2953e-05, 2.2961e-05, 2.2972e-05, 2.2983e-05, 
    2.2996e-05, 2.3007e-05, 2.3015e-05, 2.3022e-05, 2.3027e-05, 2.3027e-05, 
    2.3025e-05, 2.302e-05, 2.3012e-05, 2.3002e-05, 2.2991e-05, 2.2981e-05, 
    2.2974e-05, 2.297e-05, 2.2969e-05, 2.2969e-05, 2.2968e-05, 2.2967e-05, 
    2.2963e-05, 2.2957e-05, 2.2945e-05, 2.2931e-05, 2.2909e-05, 2.2885e-05, 
    2.2856e-05, 2.2825e-05, 2.2793e-05, 2.2761e-05, 2.2733e-05, 2.2711e-05, 
    2.2694e-05, 2.2679e-05, 2.267e-05, 2.2662e-05, 2.2658e-05, 2.2659e-05, 
    2.2662e-05, 2.267e-05, 2.2678e-05, 2.2688e-05, 2.2698e-05, 2.2708e-05, 
    2.2716e-05, 2.2723e-05, 2.2723e-05, 2.2721e-05, 2.2716e-05, 2.2709e-05, 
    2.2702e-05, 2.2694e-05, 2.2688e-05, 2.2682e-05, 2.2677e-05, 2.2673e-05, 
    2.267e-05, 2.2668e-05, 2.2667e-05, 2.2667e-05, 2.2667e-05, 2.2667e-05, 
    2.2666e-05, 2.2665e-05, 2.2664e-05, 2.2663e-05, 2.2664e-05, 2.2666e-05, 
    2.2667e-05, 2.2669e-05, 2.2671e-05, 2.2673e-05, 2.2675e-05, 2.2677e-05, 
    2.2679e-05, 2.2681e-05, 2.2686e-05, 2.2694e-05, 2.2706e-05, 2.2719e-05, 
    2.2734e-05, 2.2747e-05, 2.2759e-05, 2.2769e-05, 2.2769e-05, 2.2761e-05, 
    2.2748e-05, 2.2734e-05, 2.2716e-05, 2.2696e-05, 2.2674e-05, 2.2655e-05, 
    2.2638e-05, 2.2624e-05, 2.2611e-05, 2.2598e-05, 2.2588e-05, 2.2579e-05, 
    2.2573e-05, 2.2568e-05, 2.2564e-05, 2.2555e-05, 2.2545e-05, 2.253e-05, 
    2.251e-05, 2.2483e-05, 2.2445e-05, 2.2402e-05, 2.235e-05, 2.2295e-05, 
    2.2231e-05, 2.2159e-05, 2.2082e-05, 2.2011e-05, 2.1944e-05, 2.1887e-05, 
    2.1825e-05, 2.1761e-05, 2.1688e-05, 2.1617e-05, 2.155e-05, 2.1491e-05, 
    2.1436e-05, 2.1379e-05, 2.1318e-05, 2.1243e-05, 2.1153e-05, 2.1049e-05, 
    2.0921e-05, 2.0788e-05, 2.0649e-05, 2.0514e-05, 2.0384e-05, 2.0258e-05, 
    2.0133e-05, 2.0013e-05, 1.9889e-05, 1.9761e-05, 1.9638e-05, 1.9519e-05, 
    1.9427e-05, 1.9339e-05, 1.9259e-05, 1.9178e-05, 1.9096e-05, 1.9025e-05, 
    1.8959e-05, 1.8902e-05, 1.8847e-05, 1.8792e-05, 1.8752e-05, 1.8716e-05, 
    1.8693e-05, 1.8679e-05, 1.8672e-05, 1.8673e-05, 1.8675e-05, 1.8678e-05, 
    1.8685e-05, 1.8694e-05, 1.8707e-05, 1.8722e-05, 1.874e-05, 1.8762e-05, 
    1.8788e-05, 1.8819e-05, 1.8853e-05, 1.8893e-05, 1.893e-05, 1.8964e-05, 
    1.8991e-05, 1.9016e-05, 1.9031e-05, 1.9043e-05, 1.9048e-05, 1.9046e-05, 
    1.9042e-05, 1.903e-05, 1.9019e-05, 1.9008e-05, 1.8998e-05, 1.8988e-05, 
    1.897e-05, 1.8952e-05, 1.8933e-05, 1.8914e-05, 1.8896e-05, 1.8864e-05, 
    1.8825e-05, 1.8772e-05, 1.8725e-05, 1.8681e-05, 1.8668e-05, 1.866e-05, 
    1.8664e-05, 1.8669e-05, 1.8675e-05, 1.8677e-05, 1.8676e-05, 1.8673e-05, 
    1.8674e-05, 1.8678e-05, 1.8687e-05, 1.8697e-05, 1.8704e-05, 1.8711e-05, 
    1.8717e-05, 1.8719e-05, 1.872e-05, 1.8719e-05, 1.872e-05, 1.8723e-05, 
    1.8729e-05, 1.8736e-05, 1.8745e-05, 1.8752e-05, 1.8755e-05, 1.8755e-05, 
    1.8752e-05, 1.8746e-05, 1.8742e-05, 1.8741e-05, 1.8745e-05, 1.8752e-05, 
    1.8765e-05, 1.878e-05, 1.8797e-05, 1.8809e-05, 1.8817e-05, 1.8808e-05, 
    1.8794e-05, 1.8772e-05, 1.8745e-05, 1.8713e-05, 1.8672e-05, 1.8628e-05, 
    1.8577e-05, 1.8529e-05, 1.8484e-05, 1.8459e-05, 1.844e-05, 1.8434e-05, 
    1.843e-05, 1.8431e-05, 1.8436e-05, 1.8441e-05, 1.8448e-05, 1.8454e-05, 
    1.846e-05, 1.8464e-05, 1.8466e-05, 1.8467e-05, 1.8468e-05, 1.8467e-05, 
    1.8462e-05, 1.8456e-05, 1.8448e-05, 1.8439e-05, 1.843e-05, 1.8424e-05, 
    1.842e-05, 1.8416e-05, 1.8412e-05, 1.8409e-05, 1.8407e-05, 1.8404e-05, 
    1.8404e-05, 1.8407e-05, 1.8421e-05, 1.8444e-05, 1.8474e-05, 1.8513e-05, 
    1.8553e-05, 1.8591e-05, 1.8625e-05, 1.8656e-05, 1.8678e-05, 1.8695e-05, 
    1.87e-05, 1.8698e-05, 1.869e-05, 1.8661e-05, 1.8624e-05, 1.8571e-05, 
    1.8512e-05, 1.8446e-05, 1.8384e-05, 1.8325e-05, 1.8282e-05, 1.8244e-05, 
    1.8217e-05, 1.8203e-05, 1.8195e-05, 1.8187e-05, 1.8178e-05, 1.8168e-05, 
    1.8141e-05, 1.8104e-05, 1.8035e-05, 1.7958e-05, 1.7863e-05, 1.776e-05, 
    1.7651e-05, 1.7553e-05, 1.7461e-05, 1.7387e-05, 1.7324e-05, 1.7271e-05, 
    1.7235e-05, 1.7203e-05, 1.7175e-05, 1.7146e-05, 1.7117e-05, 1.709e-05, 
    1.7062e-05, 1.7037e-05, 1.7011e-05, 1.6985e-05, 1.6961e-05, 1.6937e-05, 
    1.6921e-05, 1.6908e-05, 1.6898e-05, 1.6892e-05, 1.6888e-05, 1.6883e-05, 
    1.6877e-05, 1.6867e-05, 1.6855e-05, 1.6841e-05, 1.6824e-05, 1.6807e-05, 
    1.6792e-05, 1.6777e-05, 1.6763e-05, 1.6742e-05, 1.6723e-05, 1.6706e-05, 
    1.6691e-05, 1.6678e-05, 1.667e-05, 1.6663e-05, 1.6657e-05, 1.6649e-05, 
    1.664e-05, 1.6627e-05, 1.6613e-05, 1.6601e-05, 1.6591e-05, 1.6584e-05, 
    1.6582e-05, 1.6583e-05, 1.6589e-05, 1.66e-05, 1.6615e-05, 1.6631e-05, 
    1.6647e-05, 1.6657e-05, 1.6664e-05, 1.6668e-05, 1.6672e-05, 1.6677e-05, 
    1.6683e-05, 1.6687e-05, 1.6688e-05, 1.6687e-05, 1.6683e-05, 1.6674e-05, 
    1.6665e-05, 1.6656e-05, 1.6648e-05, 1.6641e-05, 1.663e-05, 1.6617e-05, 
    1.6597e-05, 1.6579e-05, 1.6562e-05, 1.6548e-05, 1.6535e-05, 1.6522e-05, 
    1.651e-05, 1.6498e-05, 1.6484e-05, 1.647e-05, 1.6457e-05, 1.6446e-05, 
    1.6436e-05, 1.6427e-05, 1.6418e-05, 1.641e-05, 1.6402e-05, 1.6395e-05, 
    1.639e-05, 1.6386e-05, 1.6385e-05, 1.6384e-05, 1.6384e-05, 1.6384e-05, 
    1.6384e-05, 1.6385e-05, 1.6385e-05, 1.6385e-05, 1.6385e-05, 1.6386e-05, 
    1.6387e-05, 1.639e-05, 1.6397e-05, 1.6407e-05, 1.6419e-05, 1.6438e-05, 
    1.646e-05, 1.6488e-05, 1.6525e-05, 1.6567e-05, 1.6621e-05, 1.6677e-05, 
    1.6738e-05, 1.6801e-05, 1.6865e-05, 1.6926e-05, 1.6985e-05, 1.7037e-05, 
    1.708e-05, 1.7117e-05, 1.7144e-05, 1.7167e-05, 1.7184e-05, 1.72e-05, 
    1.7216e-05, 1.723e-05, 1.7244e-05, 1.7254e-05, 1.7263e-05, 1.7269e-05, 
    1.7273e-05, 1.7278e-05, 1.7284e-05, 1.7292e-05, 1.7304e-05, 1.7321e-05, 
    1.7341e-05, 1.7372e-05, 1.7406e-05, 1.7447e-05, 1.7483e-05, 1.7516e-05, 
    1.7532e-05, 1.7543e-05, 1.7543e-05, 1.7542e-05, 1.7541e-05, 1.7556e-05, 
    1.7581e-05, 1.7631e-05, 1.7704e-05, 1.7793e-05, 1.7905e-05, 1.8023e-05, 
    1.8156e-05, 1.8291e-05, 1.8427e-05, 1.856e-05, 1.8692e-05, 1.8826e-05, 
    1.8961e-05, 1.9097e-05, 1.9232e-05, 1.9365e-05, 1.9489e-05, 1.9608e-05, 
    1.972e-05, 1.982e-05, 1.9917e-05, 2.002e-05, 2.0129e-05, 2.0248e-05, 
    2.0385e-05, 2.0528e-05, 2.0678e-05, 2.0829e-05, 2.0983e-05, 2.1146e-05, 
    2.1312e-05, 2.1453e-05, 2.1579e-05, 2.1674e-05, 2.1741e-05, 2.1791e-05, 
    2.1805e-05, 2.1807e-05, 2.1783e-05, 2.174e-05, 2.1682e-05, 2.1605e-05, 
    2.1522e-05, 2.1431e-05, 2.1344e-05, 2.1259e-05, 2.1184e-05, 2.1111e-05, 
    2.1045e-05, 2.0982e-05, 2.0923e-05, 2.0877e-05, 2.0834e-05, 2.0798e-05, 
    2.0767e-05, 2.0742e-05, 2.0724e-05, 2.0709e-05, 2.0696e-05, 2.0681e-05, 
    2.0663e-05, 2.064e-05, 2.0616e-05, 2.0584e-05, 2.055e-05, 2.051e-05, 
    2.0465e-05, 2.0417e-05, 2.0358e-05, 2.0294e-05, 2.0219e-05, 2.014e-05, 
    2.0058e-05, 1.9989e-05, 1.9925e-05, 1.9876e-05, 1.9839e-05, 1.9812e-05, 
    1.9798e-05, 1.9786e-05, 1.9781e-05, 1.9776e-05, 1.9774e-05, 1.9772e-05, 
    1.9771e-05, 1.9769e-05, 1.9767e-05, 1.9763e-05, 1.9755e-05, 1.9746e-05, 
    1.973e-05, 1.9712e-05, 1.969e-05, 1.9665e-05, 1.9638e-05, 1.9607e-05, 
    1.9574e-05, 1.9536e-05, 1.9502e-05, 1.9471e-05, 1.9447e-05, 1.9426e-05, 
    1.9412e-05, 1.9404e-05, 1.9399e-05, 1.9397e-05, 1.9396e-05, 1.9396e-05, 
    1.9392e-05, 1.9386e-05, 1.9375e-05, 1.9363e-05, 1.9351e-05, 1.9339e-05, 
    1.9326e-05, 1.932e-05, 1.9316e-05, 1.9314e-05, 1.9315e-05, 1.9319e-05, 
    1.9326e-05, 1.9335e-05, 1.9345e-05, 1.9356e-05, 1.9368e-05, 1.9382e-05, 
    1.9397e-05, 1.9418e-05, 1.9441e-05, 1.9464e-05, 1.9487e-05, 1.9509e-05, 
    1.9534e-05, 1.9562e-05, 1.9593e-05, 1.9626e-05, 1.966e-05, 1.97e-05, 
    1.9739e-05, 1.9776e-05, 1.9807e-05, 1.9835e-05, 1.9855e-05, 1.9872e-05, 
    1.9885e-05, 1.9897e-05, 1.9908e-05, 1.9919e-05, 1.9928e-05, 1.9936e-05, 
    1.9943e-05, 1.9948e-05, 1.9948e-05, 1.9946e-05, 1.9938e-05, 1.993e-05, 
    1.9921e-05, 1.9912e-05, 1.9906e-05, 1.9911e-05, 1.9922e-05, 1.994e-05, 
    1.9965e-05, 1.9994e-05, 2.0029e-05, 2.0069e-05, 2.0115e-05, 2.017e-05, 
    2.0228e-05, 2.0289e-05, 2.0347e-05, 2.0402e-05, 2.0448e-05, 2.0491e-05, 
    2.0523e-05, 2.0553e-05, 2.0577e-05, 2.0595e-05, 2.061e-05, 2.0618e-05, 
    2.0625e-05, 2.0629e-05, 2.0631e-05, 2.0632e-05, 2.0632e-05, 2.0632e-05, 
    2.0634e-05, 2.0636e-05, 2.064e-05, 2.0645e-05, 2.0651e-05, 2.0657e-05, 
    2.0666e-05, 2.0675e-05, 2.0688e-05, 2.0702e-05, 2.0716e-05, 2.0725e-05, 
    2.0728e-05, 2.0718e-05, 2.0705e-05, 2.0687e-05, 2.0671e-05, 2.0658e-05, 
    2.0654e-05, 2.0654e-05, 2.0661e-05, 2.0667e-05, 2.067e-05, 2.0669e-05, 
    2.0665e-05, 2.0655e-05, 2.0642e-05, 2.0625e-05, 2.0603e-05, 2.0577e-05, 
    2.0542e-05, 2.0505e-05, 2.0462e-05, 2.0414e-05, 2.0363e-05, 2.0311e-05, 
    2.0257e-05, 2.0203e-05, 2.0148e-05, 2.0092e-05, 2.005e-05, 2.0013e-05, 
    1.9987e-05, 1.9967e-05, 1.9951e-05, 1.9943e-05, 1.9937e-05, 1.9934e-05, 
    1.9934e-05, 1.9936e-05, 1.9943e-05, 1.9954e-05, 1.9973e-05, 1.9995e-05, 
    2.0023e-05, 2.0061e-05, 2.0103e-05, 2.0154e-05, 2.0206e-05, 2.0259e-05, 
    2.031e-05, 2.0361e-05, 2.0409e-05, 2.0455e-05, 2.0496e-05, 2.0539e-05, 
    2.0583e-05, 2.0639e-05, 2.0699e-05, 2.0767e-05, 2.0842e-05, 2.0921e-05, 
    2.1013e-05, 2.111e-05, 2.1222e-05, 2.1344e-05, 2.1472e-05, 2.161e-05, 
    2.1751e-05, 2.1904e-05, 2.2056e-05, 2.2209e-05, 2.2338e-05, 2.2458e-05, 
    2.2552e-05, 2.2633e-05, 2.2699e-05, 2.2751e-05, 2.2798e-05, 2.2833e-05, 
    2.2867e-05, 2.2897e-05, 2.2924e-05, 2.2949e-05, 2.2972e-05, 2.2996e-05, 
    2.3019e-05, 2.3044e-05, 2.307e-05, 2.3101e-05, 2.3132e-05, 2.3165e-05, 
    2.3199e-05, 2.3234e-05, 2.3253e-05, 2.3268e-05, 2.3271e-05, 2.3269e-05, 
    2.3264e-05, 2.3259e-05, 2.3257e-05, 2.3261e-05, 2.3273e-05, 2.3293e-05, 
    2.3328e-05, 2.3368e-05, 2.3425e-05, 2.3491e-05, 2.3568e-05, 2.3653e-05, 
    2.3738e-05, 2.382e-05, 2.3895e-05, 2.3966e-05, 2.4027e-05, 2.4086e-05, 
    2.4141e-05, 2.4196e-05, 2.4249e-05, 2.4305e-05, 2.4362e-05, 2.4423e-05, 
    2.4492e-05, 2.4572e-05, 2.4666e-05, 2.4767e-05, 2.4887e-05, 2.5012e-05, 
    2.5146e-05, 2.5283e-05, 2.5421e-05, 2.5546e-05, 2.5664e-05, 2.5767e-05, 
    2.5857e-05, 2.5939e-05, 2.6003e-05, 2.606e-05, 2.6102e-05, 2.6138e-05, 
    2.6168e-05, 2.6192e-05, 2.6213e-05, 2.6229e-05, 2.624e-05, 2.6247e-05, 
    2.6244e-05, 2.6237e-05, 2.622e-05, 2.6201e-05, 2.618e-05, 2.6161e-05, 
    2.6142e-05, 2.6125e-05, 2.6111e-05, 2.6101e-05, 2.6098e-05, 2.6098e-05, 
    2.6108e-05, 2.6119e-05, 2.6131e-05, 2.6139e-05, 2.6144e-05, 2.6145e-05, 
    2.6145e-05, 2.6143e-05, 2.614e-05, 2.6137e-05, 2.6134e-05, 2.6131e-05, 
    2.6126e-05, 2.612e-05, 2.6112e-05, 2.6099e-05, 2.6084e-05, 2.6064e-05, 
    2.6039e-05, 2.6011e-05, 2.5988e-05, 2.5968e-05, 2.5959e-05, 2.5957e-05, 
    2.596e-05, 2.5967e-05, 2.5973e-05, 2.5972e-05, 2.5962e-05, 2.5942e-05, 
    2.5905e-05, 2.5864e-05, 2.5815e-05, 2.5761e-05, 2.5702e-05, 2.5638e-05, 
    2.5573e-05, 2.5513e-05, 2.5455e-05, 2.54e-05, 2.5346e-05, 2.5293e-05, 
    2.5245e-05, 2.5201e-05, 2.5161e-05, 2.5129e-05, 2.51e-05, 2.5081e-05, 
    2.5061e-05, 2.5037e-05, 2.4995e-05, 2.4943e-05, 2.4853e-05, 2.4754e-05, 
    2.4637e-05, 2.4512e-05, 2.4381e-05, 2.4238e-05, 2.4096e-05, 2.3966e-05, 
    2.3854e-05, 2.3757e-05, 2.3693e-05, 2.3641e-05, 2.3621e-05, 2.3612e-05, 
    2.3615e-05, 2.363e-05, 2.3647e-05, 2.3664e-05, 2.3678e-05, 2.3689e-05, 
    2.3695e-05, 2.3698e-05, 2.3696e-05, 2.369e-05, 2.368e-05, 2.3667e-05, 
    2.3653e-05, 2.3635e-05, 2.3617e-05, 2.3597e-05, 2.3578e-05, 2.3558e-05, 
    2.354e-05, 2.3524e-05, 2.3513e-05, 2.3508e-05, 2.3505e-05, 2.3507e-05, 
    2.3509e-05, 2.3512e-05, 2.3514e-05, 2.3516e-05, 2.3519e-05, 2.3524e-05, 
    2.3534e-05, 2.3549e-05, 2.3568e-05, 2.3593e-05, 2.3619e-05, 2.3647e-05, 
    2.3677e-05, 2.3708e-05, 2.3742e-05, 2.3776e-05, 2.3808e-05, 2.3838e-05, 
    2.3865e-05, 2.3885e-05, 2.3902e-05, 2.3914e-05, 2.3923e-05, 2.3931e-05, 
    2.3935e-05, 2.3939e-05, 2.394e-05, 2.3942e-05, 2.3942e-05, 2.3942e-05, 
    2.3942e-05, 2.3943e-05, 2.3943e-05, 2.3944e-05, 2.3945e-05, 2.3945e-05, 
    2.3944e-05, 2.3942e-05, 2.394e-05, 2.3939e-05, 2.3938e-05, 2.3938e-05, 
    2.3938e-05, 2.3938e-05, 2.3938e-05, 2.3938e-05, 2.3937e-05, 2.3935e-05, 
    2.393e-05, 2.3924e-05, 2.3916e-05, 2.3908e-05, 2.3898e-05, 2.3888e-05, 
    2.3878e-05, 2.3868e-05, 2.3856e-05, 2.3843e-05, 2.3826e-05, 2.3809e-05, 
    2.3792e-05, 2.3773e-05, 2.3753e-05, 2.3729e-05, 2.3703e-05, 2.3673e-05, 
    2.364e-05, 2.3606e-05, 2.3573e-05, 2.3539e-05, 2.3507e-05, 2.3473e-05, 
    2.3439e-05, 2.3403e-05, 2.3366e-05, 2.3325e-05, 2.3287e-05, 2.3251e-05, 
    2.322e-05, 2.3191e-05, 2.3167e-05, 2.3145e-05, 2.3125e-05, 2.3106e-05, 
    2.3089e-05, 2.3077e-05, 2.3067e-05, 2.3061e-05, 2.3057e-05, 2.3054e-05, 
    2.3052e-05, 2.3051e-05, 2.305e-05, 2.3048e-05, 2.3044e-05, 2.3038e-05, 
    2.303e-05, 2.3018e-05, 2.3002e-05, 2.2982e-05, 2.2957e-05, 2.293e-05, 
    2.2899e-05, 2.2862e-05, 2.2821e-05, 2.2771e-05, 2.2719e-05, 2.2665e-05, 
    2.2613e-05, 2.2563e-05, 2.2521e-05, 2.2483e-05, 2.2452e-05, 2.2426e-05, 
    2.2403e-05, 2.2385e-05, 2.237e-05, 2.236e-05, 2.2354e-05, 2.2351e-05, 
    2.2351e-05, 2.2351e-05, 2.2353e-05, 2.2354e-05, 2.2354e-05, 2.2352e-05, 
    2.2349e-05, 2.2345e-05, 2.2339e-05, 2.2333e-05, 2.2325e-05, 2.2316e-05, 
    2.2305e-05, 2.2293e-05, 2.2281e-05, 2.2271e-05, 2.2264e-05, 2.2263e-05, 
    2.2265e-05, 2.2271e-05, 2.2278e-05, 2.2286e-05, 2.2296e-05, 2.2306e-05, 
    2.2317e-05, 2.2335e-05, 2.2358e-05, 2.2391e-05, 2.2429e-05, 2.2481e-05, 
    2.2542e-05, 2.2608e-05, 2.2674e-05, 2.2739e-05, 2.2798e-05, 2.2856e-05, 
    2.2914e-05, 2.2967e-05, 2.3019e-05, 2.3063e-05, 2.3104e-05, 2.3141e-05, 
    2.317e-05, 2.3197e-05, 2.3214e-05, 2.3227e-05, 2.3236e-05, 2.3241e-05, 
    2.3244e-05, 2.3244e-05, 2.3244e-05, 2.3244e-05, 2.3243e-05, 2.3243e-05, 
    2.3237e-05, 2.3229e-05, 2.3215e-05, 2.3196e-05, 2.3173e-05, 2.3138e-05, 
    2.31e-05, 2.3055e-05, 2.3008e-05, 2.2959e-05, 2.2909e-05, 2.286e-05, 
    2.2814e-05, 2.2771e-05, 2.273e-05, 2.2688e-05, 2.2644e-05, 2.2592e-05, 
    2.2535e-05, 2.2473e-05, 2.2401e-05, 2.2324e-05, 2.2239e-05, 2.2144e-05, 
    2.2039e-05, 2.1922e-05, 2.1801e-05, 2.1673e-05, 2.1541e-05, 2.1404e-05, 
    2.1269e-05, 2.1137e-05, 2.1037e-05, 2.0952e-05, 2.0891e-05, 2.0855e-05, 
    2.083e-05, 2.083e-05, 2.0836e-05, 2.0853e-05, 2.0876e-05, 2.0901e-05, 
    2.0934e-05, 2.0967e-05, 2.1e-05, 2.1026e-05, 2.1049e-05, 2.1059e-05, 
    2.1064e-05, 2.1058e-05, 2.1045e-05, 2.1028e-05, 2.1002e-05, 2.0978e-05, 
    2.0961e-05, 2.095e-05, 2.0945e-05, 2.0944e-05, 2.0945e-05, 2.0945e-05, 
    2.0941e-05, 2.0932e-05, 2.0911e-05, 2.0884e-05, 2.0841e-05, 2.079e-05, 
    2.0728e-05, 2.065e-05, 2.0568e-05, 2.0476e-05, 2.0388e-05, 2.0306e-05, 
    2.0236e-05, 2.0172e-05, 2.0124e-05, 2.008e-05, 2.0041e-05, 2.0003e-05, 
    1.9967e-05, 1.9925e-05, 1.988e-05, 1.9827e-05, 1.9758e-05, 1.9677e-05, 
    1.9566e-05, 1.9444e-05, 1.9297e-05, 1.9135e-05, 1.8961e-05, 1.8777e-05, 
    1.8594e-05, 1.8422e-05, 1.8264e-05, 1.8117e-05, 1.7993e-05, 1.7876e-05, 
    1.778e-05, 1.7696e-05, 1.7624e-05, 1.7564e-05, 1.7508e-05, 1.7456e-05, 
    1.7405e-05, 1.7357e-05, 1.7312e-05, 1.7267e-05, 1.7229e-05, 1.7194e-05, 
    1.7164e-05, 1.7136e-05, 1.7107e-05, 1.7072e-05, 1.7034e-05, 1.6992e-05, 
    1.6947e-05, 1.6901e-05, 1.685e-05, 1.6798e-05, 1.6742e-05, 1.669e-05, 
    1.6641e-05, 1.6609e-05, 1.6581e-05, 1.6564e-05, 1.6553e-05, 1.6548e-05, 
    1.6551e-05, 1.6555e-05, 1.6562e-05, 1.657e-05, 1.6579e-05, 1.6591e-05, 
    1.6604e-05, 1.662e-05, 1.6641e-05, 1.6666e-05, 1.6699e-05, 1.6736e-05, 
    1.6781e-05, 1.6828e-05, 1.6879e-05, 1.6928e-05, 1.6977e-05, 1.7022e-05, 
    1.7067e-05, 1.7111e-05, 1.715e-05, 1.7186e-05, 1.7204e-05, 1.7215e-05, 
    1.7214e-05, 1.7202e-05, 1.7185e-05, 1.7152e-05, 1.7114e-05, 1.7062e-05, 
    1.6999e-05, 1.6929e-05, 1.6856e-05, 1.6783e-05, 1.6717e-05, 1.6659e-05, 
    1.6606e-05, 1.6568e-05, 1.6535e-05, 1.6517e-05, 1.6508e-05, 1.6509e-05, 
    1.6533e-05, 1.6566e-05, 1.6622e-05, 1.6685e-05, 1.6758e-05, 1.6827e-05, 
    1.689e-05, 1.6925e-05, 1.6949e-05, 1.696e-05, 1.6963e-05, 1.6961e-05, 
    1.6954e-05, 1.6943e-05, 1.6927e-05, 1.6905e-05, 1.6882e-05, 1.6861e-05, 
    1.6844e-05, 1.6834e-05, 1.6831e-05, 1.6833e-05, 1.6844e-05, 1.6856e-05, 
    5.2279e-06, 5.2153e-06, 5.1993e-06, 5.1802e-06, 5.1583e-06, 5.1335e-06, 
    5.1063e-06, 5.0769e-06, 5.0454e-06, 5.0123e-06, 4.9776e-06, 4.9418e-06, 
    4.9049e-06, 4.8673e-06, 4.8293e-06, 4.791e-06, 4.7528e-06, 4.7149e-06, 
    4.6774e-06, 4.6407e-06, 4.605e-06, 4.5704e-06, 4.5371e-06, 4.5054e-06, 
    4.4754e-06, 4.4472e-06, 4.4209e-06, 4.3968e-06, 4.3749e-06, 4.3553e-06, 
    4.3382e-06, 4.3235e-06, 4.3114e-06, 4.302e-06, 4.2954e-06, 4.2916e-06, 
    4.2907e-06, 4.2928e-06, 4.2979e-06, 4.3063e-06, 4.3176e-06, 4.3325e-06, 
    4.3506e-06, 4.3721e-06, 4.3971e-06, 4.4256e-06, 4.4576e-06, 4.493e-06, 
    4.532e-06, 4.5742e-06, 4.6196e-06, 4.668e-06, 4.7191e-06, 4.7725e-06, 
    4.8281e-06, 4.8852e-06, 4.9433e-06, 5.0019e-06, 5.0602e-06, 5.1175e-06, 
    5.1732e-06, 5.2263e-06, 5.2761e-06, 5.3216e-06, 5.3623e-06, 5.3972e-06, 
    5.4259e-06, 5.4475e-06, 5.4617e-06, 5.4681e-06, 5.4663e-06, 5.4564e-06, 
    5.4383e-06, 5.4125e-06, 5.3789e-06, 5.3385e-06, 5.2918e-06, 5.2393e-06, 
    5.1821e-06, 5.1211e-06, 5.0572e-06, 4.9915e-06, 4.9248e-06, 4.8582e-06, 
    4.7926e-06, 4.7289e-06, 4.6679e-06, 4.6103e-06, 4.5567e-06, 4.5076e-06, 
    4.4635e-06, 4.4248e-06, 4.3918e-06, 4.3645e-06, 4.3432e-06, 4.3279e-06, 
    4.3185e-06, 4.315e-06, 4.3171e-06, 4.3247e-06, 4.3375e-06, 4.3552e-06, 
    4.3773e-06, 4.4035e-06, 4.4332e-06, 4.4661e-06, 4.5015e-06, 4.5388e-06, 
    4.5775e-06, 4.6169e-06, 4.6564e-06, 4.6955e-06, 4.7334e-06, 4.7696e-06, 
    4.8035e-06, 4.8346e-06, 4.8624e-06, 4.8866e-06, 4.9069e-06, 4.9229e-06, 
    4.9347e-06, 4.9421e-06, 4.945e-06, 4.9436e-06, 4.9381e-06, 4.9288e-06, 
    4.9158e-06, 4.8996e-06, 4.8806e-06, 4.859e-06, 4.8354e-06, 4.81e-06, 
    4.7834e-06, 4.7557e-06, 4.7275e-06, 4.6988e-06, 4.6701e-06, 4.6413e-06, 
    4.6129e-06, 4.5848e-06, 4.5572e-06, 4.5301e-06, 4.5035e-06, 4.4773e-06, 
    4.4516e-06, 4.4263e-06, 4.4015e-06, 4.3771e-06, 4.3529e-06, 4.329e-06, 
    4.3055e-06, 4.2823e-06, 4.2595e-06, 4.2371e-06, 4.2151e-06, 4.1936e-06, 
    4.1728e-06, 4.1527e-06, 4.1334e-06, 4.1149e-06, 4.0973e-06, 4.0807e-06, 
    4.0652e-06, 4.0508e-06, 4.0375e-06, 4.0253e-06, 4.0142e-06, 4.0043e-06, 
    3.9954e-06, 3.9877e-06, 3.9809e-06, 3.975e-06, 3.9701e-06, 3.966e-06, 
    3.9626e-06, 3.9599e-06, 3.9578e-06, 3.9562e-06, 3.955e-06, 3.9543e-06, 
    3.9538e-06, 3.9535e-06, 3.9534e-06, 3.9534e-06, 3.9533e-06, 3.9533e-06, 
    3.953e-06, 3.9525e-06, 3.9515e-06, 3.9501e-06, 3.9482e-06, 3.9454e-06, 
    3.9418e-06, 3.9371e-06, 3.9315e-06, 3.9245e-06, 3.9163e-06, 3.9067e-06, 
    3.8957e-06, 3.8833e-06, 3.8694e-06, 3.8542e-06, 3.8376e-06, 3.8198e-06, 
    3.801e-06, 3.7812e-06, 3.7605e-06, 3.7392e-06, 3.7173e-06, 3.6949e-06, 
    3.6724e-06, 3.6496e-06, 3.6267e-06, 3.6038e-06, 3.581e-06, 3.5583e-06, 
    3.5357e-06, 3.5134e-06, 3.4914e-06, 3.4697e-06, 3.4483e-06, 3.4274e-06, 
    3.407e-06, 3.3872e-06, 3.3681e-06, 3.3498e-06, 3.3324e-06, 3.3161e-06, 
    3.3009e-06, 3.287e-06, 3.2745e-06, 3.2635e-06, 3.2541e-06, 3.2465e-06, 
    3.2406e-06, 3.2365e-06, 3.2343e-06, 3.234e-06, 3.2356e-06, 3.2391e-06, 
    3.2445e-06, 3.2516e-06, 3.2605e-06, 3.2711e-06, 3.2831e-06, 3.2966e-06, 
    3.3115e-06, 3.3275e-06, 3.3446e-06, 3.3626e-06, 3.3814e-06, 3.4008e-06, 
    3.4208e-06, 3.4413e-06, 3.4621e-06, 3.4832e-06, 3.5046e-06, 3.5262e-06, 
    3.548e-06, 3.57e-06, 3.5922e-06, 3.6147e-06, 3.6374e-06, 3.6604e-06, 
    3.6837e-06, 3.7074e-06, 3.7313e-06, 3.7556e-06, 3.78e-06, 3.8046e-06, 
    3.8292e-06, 3.8536e-06, 3.8776e-06, 3.901e-06, 3.9236e-06, 3.945e-06, 
    3.9648e-06, 3.983e-06, 3.9989e-06, 4.0126e-06, 4.0234e-06, 4.0314e-06, 
    4.0361e-06, 4.0374e-06, 4.0353e-06, 4.0296e-06, 4.0204e-06, 4.0077e-06, 
    3.9917e-06, 3.9725e-06, 3.9504e-06, 3.9257e-06, 3.8987e-06, 3.8698e-06, 
    3.8393e-06, 3.8077e-06, 3.775e-06, 3.742e-06, 3.7086e-06, 3.6754e-06, 
    3.6425e-06, 3.6101e-06, 3.5783e-06, 3.5474e-06, 3.5174e-06, 3.4883e-06, 
    3.4602e-06, 3.4331e-06, 3.4069e-06, 3.3816e-06, 3.3574e-06, 3.3339e-06, 
    3.3113e-06, 3.2896e-06, 3.2685e-06, 3.2483e-06, 3.2287e-06, 3.2099e-06, 
    3.1918e-06, 3.1743e-06, 3.1577e-06, 3.1416e-06, 3.1263e-06, 3.1117e-06, 
    3.0978e-06, 3.0846e-06, 3.0721e-06, 3.0604e-06, 3.0494e-06, 3.0391e-06, 
    3.0295e-06, 3.0208e-06, 3.0129e-06, 3.0058e-06, 2.9996e-06, 2.9943e-06, 
    2.9899e-06, 2.9865e-06, 2.9841e-06, 2.9827e-06, 2.9823e-06, 2.9828e-06, 
    2.9843e-06, 2.9868e-06, 2.9901e-06, 2.9943e-06, 2.9992e-06, 3.0049e-06, 
    3.0111e-06, 3.0178e-06, 3.025e-06, 3.0325e-06, 3.0403e-06, 3.0483e-06, 
    3.0565e-06, 3.0647e-06, 3.0729e-06, 3.0812e-06, 3.0893e-06, 3.0973e-06, 
    3.1053e-06, 3.1131e-06, 3.1207e-06, 3.1283e-06, 3.1356e-06, 3.1428e-06, 
    3.1499e-06, 3.1568e-06, 3.1636e-06, 3.1703e-06, 3.1769e-06, 3.1835e-06, 
    3.1902e-06, 3.1969e-06, 3.2038e-06, 3.2108e-06, 3.2181e-06, 3.2257e-06, 
    3.2337e-06, 3.2421e-06, 3.251e-06, 3.2604e-06, 3.2703e-06, 3.2806e-06, 
    3.2914e-06, 3.3025e-06, 3.3139e-06, 3.3255e-06, 3.3371e-06, 3.3485e-06, 
    3.3595e-06, 3.3699e-06, 3.3795e-06, 3.3879e-06, 3.3951e-06, 3.4006e-06, 
    3.4044e-06, 3.4062e-06, 3.4058e-06, 3.4031e-06, 3.398e-06, 3.3904e-06, 
    3.3805e-06, 3.3682e-06, 3.3536e-06, 3.3369e-06, 3.3184e-06, 3.2981e-06, 
    3.2765e-06, 3.2537e-06, 3.2301e-06, 3.206e-06, 3.1816e-06, 3.1573e-06, 
    3.1333e-06, 3.1098e-06, 3.087e-06, 3.0652e-06, 3.0446e-06, 3.0252e-06, 
    3.0071e-06, 2.9904e-06, 2.9752e-06, 2.9614e-06, 2.949e-06, 2.9381e-06, 
    2.9284e-06, 2.9201e-06, 2.9129e-06, 2.9067e-06, 2.9015e-06, 2.8971e-06, 
    2.8934e-06, 2.8902e-06, 2.8875e-06, 2.8851e-06, 2.883e-06, 2.8809e-06, 
    2.879e-06, 2.877e-06, 2.8749e-06, 2.8728e-06, 2.8706e-06, 2.8682e-06, 
    2.8658e-06, 2.8634e-06, 2.8611e-06, 2.8587e-06, 2.8565e-06, 2.8545e-06, 
    2.8527e-06, 2.8513e-06, 2.8501e-06, 2.8492e-06, 2.8486e-06, 2.8483e-06, 
    2.8482e-06, 2.8483e-06, 2.8483e-06, 2.8483e-06, 2.8482e-06, 2.8476e-06, 
    2.8466e-06, 2.845e-06, 2.8427e-06, 2.8395e-06, 2.8353e-06, 2.83e-06, 
    2.8237e-06, 2.8162e-06, 2.8076e-06, 2.798e-06, 2.7874e-06, 2.7759e-06, 
    2.7639e-06, 2.7512e-06, 2.7383e-06, 2.7254e-06, 2.7125e-06, 2.7001e-06, 
    2.6883e-06, 2.6774e-06, 2.6676e-06, 2.659e-06, 2.6519e-06, 2.6464e-06, 
    2.6426e-06, 2.6406e-06, 2.6405e-06, 2.6423e-06, 2.646e-06, 2.6515e-06, 
    2.6588e-06, 2.6678e-06, 2.6782e-06, 2.6898e-06, 2.7026e-06, 2.7162e-06, 
    2.7303e-06, 2.7447e-06, 2.7591e-06, 2.773e-06, 2.7864e-06, 2.7988e-06, 
    2.81e-06, 2.8198e-06, 2.8279e-06, 2.8341e-06, 2.8384e-06, 2.8407e-06, 
    2.841e-06, 2.839e-06, 2.8351e-06, 2.8293e-06, 2.8216e-06, 2.8121e-06, 
    2.8012e-06, 2.7888e-06, 2.7751e-06, 2.7604e-06, 2.7448e-06, 2.7285e-06, 
    2.7115e-06, 2.6942e-06, 2.6765e-06, 2.6587e-06, 2.6408e-06, 2.623e-06, 
    2.6055e-06, 2.5882e-06, 2.5714e-06, 2.5552e-06, 2.5395e-06, 2.5247e-06, 
    2.5107e-06, 2.4976e-06, 2.4856e-06, 2.4748e-06, 2.4651e-06, 2.4567e-06, 
    2.4496e-06, 2.4438e-06, 2.4394e-06, 2.4364e-06, 2.4346e-06, 2.4342e-06, 
    2.435e-06, 2.437e-06, 2.4399e-06, 2.4439e-06, 2.4487e-06, 2.4542e-06, 
    2.4602e-06, 2.4667e-06, 2.4735e-06, 2.4804e-06, 2.4875e-06, 2.4946e-06, 
    2.5017e-06, 2.5086e-06, 2.5153e-06, 2.522e-06, 2.5285e-06, 2.5348e-06, 
    2.5412e-06, 2.5475e-06, 2.5539e-06, 2.5605e-06, 2.5673e-06, 2.5743e-06, 
    2.5816e-06, 2.5892e-06, 2.5971e-06, 2.6054e-06, 2.6139e-06, 2.6226e-06, 
    2.6313e-06, 2.64e-06, 2.6486e-06, 2.6568e-06, 2.6644e-06, 2.6714e-06, 
    2.6774e-06, 2.6823e-06, 2.6858e-06, 2.6878e-06, 2.6881e-06, 2.6865e-06, 
    2.683e-06, 2.6775e-06, 2.6699e-06, 2.6602e-06, 2.6486e-06, 2.6351e-06, 
    2.6199e-06, 2.603e-06, 2.5849e-06, 2.5658e-06, 2.5458e-06, 2.5254e-06, 
    2.5049e-06, 2.4844e-06, 2.4644e-06, 2.445e-06, 2.4266e-06, 2.4094e-06, 
    2.3936e-06, 2.3792e-06, 2.3665e-06, 2.3556e-06, 2.3464e-06, 2.339e-06, 
    2.3333e-06, 2.3294e-06, 2.327e-06, 2.3262e-06, 2.3266e-06, 2.3283e-06, 
    2.3311e-06, 2.3346e-06, 2.3387e-06, 2.3433e-06, 2.348e-06, 2.3528e-06, 
    2.3575e-06, 2.3618e-06, 2.3657e-06, 2.369e-06, 2.3716e-06, 2.3734e-06, 
    2.3745e-06, 2.3749e-06, 2.3744e-06, 2.3733e-06, 2.3715e-06, 2.3692e-06, 
    2.3664e-06, 2.3633e-06, 2.3599e-06, 2.3565e-06, 2.3531e-06, 2.3498e-06, 
    2.3468e-06, 2.3443e-06, 2.3422e-06, 2.3406e-06, 2.3397e-06, 2.3395e-06, 
    2.34e-06, 2.3412e-06, 2.3433e-06, 2.346e-06, 2.3496e-06, 2.3538e-06, 
    2.3586e-06, 2.3641e-06, 2.37e-06, 2.3764e-06, 2.3831e-06, 2.39e-06, 
    2.3971e-06, 2.4041e-06, 2.411e-06, 2.4176e-06, 2.4239e-06, 2.4297e-06, 
    2.4349e-06, 2.4394e-06, 2.4431e-06, 2.446e-06, 2.448e-06, 2.449e-06, 
    2.449e-06, 2.448e-06, 2.4459e-06, 2.4428e-06, 2.4388e-06, 2.4337e-06, 
    2.4277e-06, 2.4208e-06, 2.413e-06, 2.4044e-06, 2.3949e-06, 2.3848e-06, 
    2.3739e-06, 2.3624e-06, 2.3504e-06, 2.3379e-06, 2.3249e-06, 2.3115e-06, 
    2.2979e-06, 2.284e-06, 2.2701e-06, 2.2562e-06, 2.2424e-06, 2.2288e-06, 
    2.2155e-06, 2.2027e-06, 2.1903e-06, 2.1787e-06, 2.1677e-06, 2.1576e-06, 
    2.1485e-06, 2.1404e-06, 2.1333e-06, 2.1274e-06, 2.1227e-06, 2.1191e-06, 
    2.1168e-06, 2.1158e-06, 2.1159e-06, 2.1172e-06, 2.1197e-06, 2.1232e-06, 
    2.1276e-06, 2.133e-06, 2.1392e-06, 2.1459e-06, 2.1532e-06, 2.161e-06, 
    2.1689e-06, 2.1769e-06, 2.1848e-06, 2.1926e-06, 2.2e-06, 2.207e-06, 
    2.2134e-06, 2.2192e-06, 2.2244e-06, 2.2288e-06, 2.2325e-06, 2.2354e-06, 
    2.2377e-06, 2.2393e-06, 2.2403e-06, 2.2406e-06, 2.2405e-06, 2.2399e-06, 
    2.2389e-06, 2.2375e-06, 2.2358e-06, 2.2338e-06, 2.2316e-06, 2.2292e-06, 
    2.2265e-06, 2.2238e-06, 2.2209e-06, 2.2178e-06, 2.2146e-06, 2.2114e-06, 
    2.2081e-06, 2.2049e-06, 2.2017e-06, 2.1986e-06, 2.1957e-06, 2.1931e-06, 
    2.1908e-06, 2.1888e-06, 2.1873e-06, 2.1862e-06, 2.1857e-06, 2.1858e-06, 
    2.1864e-06, 2.1877e-06, 2.1895e-06, 2.1918e-06, 2.1947e-06, 2.198e-06, 
    2.2017e-06, 2.2057e-06, 2.2098e-06, 2.214e-06, 2.2181e-06, 2.222e-06, 
    2.2256e-06, 2.2287e-06, 2.2311e-06, 2.2329e-06, 2.2338e-06, 2.2339e-06, 
    2.233e-06, 2.2311e-06, 2.2281e-06, 2.2242e-06, 2.2192e-06, 2.2134e-06, 
    2.2067e-06, 2.1993e-06, 2.1912e-06, 2.1826e-06, 2.1736e-06, 2.1644e-06, 
    2.155e-06, 2.1457e-06, 2.1365e-06, 2.1275e-06, 2.119e-06, 2.111e-06, 
    2.1035e-06, 2.0966e-06, 2.0905e-06, 2.0851e-06, 2.0804e-06, 2.0766e-06, 
    2.0735e-06, 2.0713e-06, 2.0697e-06, 2.0688e-06, 2.0686e-06, 2.0689e-06, 
    2.0697e-06, 2.0709e-06, 2.0724e-06, 2.0741e-06, 2.0759e-06, 2.0778e-06, 
    2.0796e-06, 2.0813e-06, 2.0827e-06, 2.0839e-06, 2.0848e-06, 2.0853e-06, 
    2.0855e-06, 2.0853e-06, 2.0848e-06, 2.0839e-06, 2.0828e-06, 2.0814e-06, 
    2.0798e-06, 2.0781e-06, 2.0762e-06, 2.0743e-06, 2.0725e-06, 2.0706e-06, 
    2.0688e-06, 2.0671e-06, 2.0655e-06, 2.0641e-06, 2.0627e-06, 2.0615e-06, 
    2.0604e-06, 2.0594e-06, 2.0585e-06, 2.0576e-06, 2.0569e-06, 2.0562e-06, 
    2.0555e-06, 2.0548e-06, 2.0542e-06, 2.0537e-06, 2.0531e-06, 2.0526e-06, 
    2.0521e-06, 2.0516e-06, 2.0512e-06, 2.0508e-06, 2.0504e-06, 2.05e-06, 
    2.0497e-06, 2.0493e-06, 2.0489e-06, 2.0486e-06, 2.0481e-06, 2.0477e-06, 
    2.0471e-06, 2.0465e-06, 2.0458e-06, 2.045e-06, 2.0441e-06, 2.0431e-06, 
    2.0421e-06, 2.0409e-06, 2.0396e-06, 2.0383e-06, 2.0369e-06, 2.0355e-06, 
    2.0341e-06, 2.0326e-06, 2.0312e-06, 2.0298e-06, 2.0284e-06, 2.027e-06, 
    2.0257e-06, 2.0245e-06, 2.0233e-06, 2.0222e-06, 2.0211e-06, 2.0202e-06, 
    2.0193e-06, 2.0185e-06, 2.0178e-06, 2.0172e-06, 2.0168e-06, 2.0165e-06, 
    2.0163e-06, 2.0164e-06, 2.0166e-06, 2.017e-06, 2.0177e-06, 2.0186e-06, 
    2.0198e-06, 2.0212e-06, 2.0229e-06, 2.0248e-06, 2.0269e-06, 2.0292e-06, 
    2.0317e-06, 2.0343e-06, 2.037e-06, 2.0397e-06, 2.0423e-06, 2.0449e-06, 
    2.0474e-06, 2.0496e-06, 2.0516e-06, 2.0533e-06, 2.0546e-06, 2.0555e-06, 
    2.0561e-06, 2.0562e-06, 2.0559e-06, 2.0552e-06, 2.0542e-06, 2.0527e-06, 
    2.0509e-06, 2.0488e-06, 2.0465e-06, 2.044e-06, 2.0414e-06, 2.0386e-06, 
    2.036e-06, 2.0333e-06, 2.0308e-06, 2.0284e-06, 2.0262e-06, 2.0242e-06, 
    2.0225e-06, 2.0211e-06, 2.0199e-06, 2.019e-06, 2.0185e-06, 2.0182e-06, 
    2.0181e-06, 2.0183e-06, 2.0187e-06, 2.0192e-06, 2.0199e-06, 2.0207e-06, 
    2.0215e-06, 2.0224e-06, 2.0233e-06, 2.0241e-06, 2.025e-06, 2.0257e-06, 
    2.0264e-06, 2.0271e-06, 2.0276e-06, 2.0281e-06, 2.0285e-06, 2.0289e-06, 
    2.0292e-06, 2.0295e-06, 2.0297e-06, 2.0299e-06, 2.0301e-06, 2.0303e-06, 
    2.0304e-06, 2.0305e-06, 2.0306e-06, 2.0306e-06, 2.0306e-06, 2.0305e-06, 
    2.0304e-06, 2.0302e-06, 2.0299e-06, 2.0295e-06, 2.029e-06, 2.0284e-06, 
    2.0277e-06, 2.0269e-06, 2.026e-06, 2.0251e-06, 2.0241e-06, 2.0229e-06, 
    2.0218e-06, 2.0207e-06, 2.0195e-06, 2.0183e-06, 2.0171e-06, 2.0159e-06, 
    2.0147e-06, 2.0136e-06, 2.0124e-06, 2.0113e-06, 2.0102e-06, 2.009e-06, 
    2.0079e-06, 2.0068e-06, 2.0056e-06, 2.0045e-06, 2.0032e-06, 2.002e-06, 
    2.0006e-06, 1.9992e-06, 1.9977e-06, 1.9962e-06, 1.9945e-06, 1.9928e-06, 
    1.991e-06, 1.989e-06, 1.987e-06, 1.9849e-06, 1.9826e-06, 1.9803e-06, 
    1.9779e-06, 1.9754e-06, 1.9728e-06, 1.9701e-06, 1.9675e-06, 1.9647e-06, 
    1.962e-06, 1.9593e-06, 1.9567e-06, 1.9541e-06, 1.9517e-06, 1.9494e-06, 
    1.9472e-06, 1.9453e-06, 1.9436e-06, 1.9421e-06, 1.9409e-06, 1.94e-06, 
    1.9393e-06, 1.939e-06, 1.939e-06, 1.9393e-06, 1.9399e-06, 1.9408e-06, 
    1.9419e-06, 1.9433e-06, 1.9448e-06, 1.9466e-06, 1.9484e-06, 1.9504e-06, 
    1.9525e-06, 1.9547e-06, 1.9569e-06, 1.9591e-06, 1.9612e-06, 1.9634e-06, 
    1.9654e-06, 1.9674e-06, 1.9693e-06, 1.9712e-06, 1.9729e-06, 1.9745e-06, 
    1.9759e-06, 1.9773e-06, 1.9785e-06, 1.9796e-06, 1.9806e-06, 1.9815e-06, 
    1.9823e-06, 1.9829e-06, 1.9834e-06, 1.9839e-06, 1.9842e-06, 1.9844e-06, 
    1.9846e-06, 1.9846e-06, 1.9846e-06, 1.9844e-06, 1.9843e-06, 1.984e-06, 
    1.9837e-06, 1.9833e-06, 1.9828e-06, 1.9823e-06, 1.9818e-06, 1.9812e-06, 
    1.9806e-06, 1.9799e-06, 1.9792e-06, 1.9784e-06, 1.9776e-06, 1.9768e-06, 
    1.9759e-06, 1.975e-06, 1.974e-06, 1.973e-06, 1.9719e-06, 1.9708e-06, 
    1.9696e-06, 1.9683e-06, 1.967e-06, 1.9656e-06, 1.9641e-06, 1.9625e-06, 
    1.9609e-06, 1.9592e-06, 1.9575e-06, 1.9558e-06, 1.954e-06, 1.9523e-06, 
    1.9506e-06, 1.9488e-06, 1.9472e-06, 1.9456e-06, 1.944e-06, 1.9426e-06, 
    1.9412e-06, 1.94e-06, 1.9389e-06, 1.9378e-06, 1.9369e-06, 1.9361e-06, 
    1.9355e-06, 1.9349e-06, 1.9344e-06, 1.9341e-06, 1.9339e-06, 1.9338e-06, 
    1.9338e-06, 1.9339e-06, 1.9341e-06, 1.9344e-06, 1.9349e-06, 1.9354e-06, 
    1.9361e-06, 1.9369e-06, 1.9377e-06, 1.9387e-06, 1.9396e-06, 1.9407e-06, 
    1.9419e-06, 1.943e-06, 1.9441e-06, 1.9452e-06, 1.9463e-06, 1.9473e-06, 
    1.9482e-06, 1.949e-06, 1.9496e-06, 1.95e-06, 1.9503e-06, 1.9504e-06, 
    1.9503e-06, 1.95e-06, 1.9496e-06, 1.9489e-06, 1.9481e-06, 1.9472e-06, 
    1.9461e-06, 1.945e-06, 1.9438e-06, 1.9425e-06, 1.9413e-06, 1.94e-06, 
    1.9389e-06, 1.9377e-06, 1.9367e-06, 1.9358e-06, 1.9349e-06, 1.9342e-06, 
    1.9336e-06, 1.9332e-06, 1.9329e-06, 1.9326e-06, 1.9325e-06, 1.9325e-06, 
    1.9326e-06, 1.9328e-06, 1.933e-06, 1.9332e-06, 1.9336e-06, 1.9339e-06, 
    1.9343e-06, 1.9347e-06, 1.9351e-06, 1.9354e-06, 1.9358e-06, 1.9362e-06, 
    1.9365e-06, 1.9369e-06, 1.9372e-06, 1.9375e-06, 1.9378e-06, 1.938e-06, 
    1.9382e-06, 1.9382e-06, 1.9383e-06, 1.9383e-06, 1.9381e-06, 1.9379e-06, 
    1.9376e-06, 1.9371e-06, 1.9365e-06, 1.9357e-06, 1.9348e-06, 1.9338e-06, 
    1.9326e-06, 1.9314e-06, 1.9301e-06, 1.9288e-06, 1.9275e-06, 1.9263e-06, 
    1.9253e-06, 1.9244e-06, 1.9239e-06, 1.9236e-06, 1.9238e-06, 1.9244e-06, 
    1.9255e-06, 1.9271e-06, 1.9292e-06, 1.9319e-06, 1.9351e-06, 1.9388e-06, 
    1.943e-06, 1.9475e-06, 1.9523e-06, 1.9573e-06, 1.9623e-06, 1.9673e-06, 
    1.9721e-06, 1.9765e-06, 1.9805e-06, 1.9839e-06, 1.9867e-06, 1.9886e-06, 
    1.9897e-06, 1.99e-06, 1.9893e-06, 1.9877e-06, 1.9853e-06, 1.982e-06, 
    1.978e-06, 1.9734e-06, 1.9682e-06, 1.9625e-06, 1.9566e-06, 1.9505e-06, 
    1.9443e-06, 1.9382e-06, 1.9323e-06, 1.9266e-06, 1.9212e-06, 1.9163e-06, 
    1.9118e-06, 1.9078e-06, 1.9043e-06, 1.9014e-06, 1.899e-06, 1.8972e-06, 
    1.8959e-06, 1.8951e-06, 1.8948e-06, 1.8949e-06, 1.8955e-06, 1.8964e-06, 
    1.8978e-06, 1.8995e-06, 1.9014e-06, 1.9037e-06, 1.9062e-06, 1.9089e-06, 
    1.9118e-06, 1.9149e-06, 1.9181e-06, 1.9214e-06, 1.9248e-06, 1.9282e-06, 
    1.9317e-06, 1.9352e-06, 1.9386e-06, 1.942e-06, 1.9452e-06, 1.9484e-06, 
    1.9514e-06, 1.9542e-06, 1.9569e-06, 1.9593e-06, 1.9616e-06, 1.9635e-06, 
    1.9653e-06, 1.9667e-06, 1.9679e-06, 1.9688e-06, 1.9695e-06, 1.9699e-06, 
    1.97e-06, 1.9699e-06, 1.9695e-06, 1.9689e-06, 1.9681e-06, 1.9671e-06, 
    1.9659e-06, 1.9645e-06, 1.9629e-06, 1.9612e-06, 1.9593e-06, 1.9573e-06, 
    1.9552e-06, 1.9528e-06, 1.9504e-06, 1.9479e-06, 1.9453e-06, 1.9425e-06, 
    1.9397e-06, 1.9368e-06, 1.9338e-06, 1.9307e-06, 1.9275e-06, 1.9242e-06, 
    1.9209e-06, 1.9176e-06, 1.9141e-06, 1.9107e-06, 1.9071e-06, 1.9036e-06, 
    1.9001e-06, 1.8966e-06, 1.8932e-06, 1.8898e-06, 1.8865e-06, 1.8834e-06, 
    1.8804e-06, 1.8775e-06, 1.8749e-06, 1.8725e-06, 1.8704e-06, 1.8685e-06, 
    1.8669e-06, 1.8656e-06, 1.8646e-06, 1.8638e-06, 1.8634e-06, 1.8633e-06, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_L1_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_L2_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 bangle_qual =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100 ;

 bangle_opt_qual =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100 ;

 alt_refrac =
  30.994, 32.49, 33.938, 35.333, 36.697, 38.061, 39.442, 40.858, 42.299, 
    43.766, 45.29, 46.898, 48.599, 50.4, 52.31, 54.349, 56.535, 58.845, 
    61.284, 63.845, 66.534, 69.355, 72.283, 75.308, 78.361, 81.447, 84.575, 
    87.755, 90.991, 94.254, 97.541, 100.85, 104.19, 107.59, 111.04, 114.56, 
    118.15, 121.81, 125.53, 129.29, 133.09, 136.92, 140.79, 144.71, 148.65, 
    152.61, 156.56, 160.49, 164.4, 168.31, 172.21, 176.1, 179.98, 183.85, 
    187.71, 191.54, 195.36, 199.15, 202.92, 206.69, 210.48, 214.29, 218.13, 
    222.01, 225.9, 229.78, 233.65, 237.51, 241.36, 245.22, 249.07, 252.92, 
    256.74, 260.53, 264.29, 268.01, 271.71, 275.41, 279.09, 282.77, 286.44, 
    290.08, 293.69, 297.31, 300.94, 304.61, 308.29, 311.98, 315.68, 319.4, 
    323.12, 326.85, 330.6, 334.37, 338.17, 341.98, 345.81, 349.64, 353.49, 
    357.35, 361.21, 365.08, 368.96, 372.83, 376.72, 380.61, 384.52, 388.43, 
    392.35, 396.27, 400.19, 404.11, 408.04, 411.97, 415.92, 419.86, 423.81, 
    427.75, 431.69, 435.61, 439.52, 443.42, 447.29, 451.15, 455.01, 458.85, 
    462.68, 466.5, 470.31, 474.12, 477.92, 481.73, 485.52, 489.32, 493.11, 
    496.91, 500.72, 504.53, 508.35, 512.18, 516.01, 519.84, 523.66, 527.49, 
    531.33, 535.16, 538.99, 542.82, 546.65, 550.48, 554.32, 558.15, 561.98, 
    565.8, 569.62, 573.47, 577.33, 581.19, 585.06, 588.95, 592.87, 596.82, 
    600.8, 604.81, 608.83, 612.88, 616.95, 621.05, 625.16, 629.29, 633.46, 
    637.65, 641.86, 646.1, 650.35, 654.62, 658.9, 663.21, 667.55, 671.92, 
    676.34, 680.79, 685.28, 689.83, 694.43, 699.12, 703.9, 708.76, 713.71, 
    718.76, 723.92, 729.19, 734.53, 739.9, 745.28, 750.65, 756.03, 761.4, 
    766.75, 772.06, 777.33, 782.55, 787.77, 793.01, 798.24, 803.48, 808.73, 
    813.99, 819.27, 824.53, 829.78, 835.02, 840.27, 845.53, 850.77, 855.96, 
    861.06, 866.11, 871.12, 876.08, 881.01, 885.9, 890.72, 895.49, 900.16, 
    904.73, 909.2, 913.56, 917.79, 921.95, 926.03, 930.05, 934.05, 938.05, 
    942.07, 946.11, 950.17, 954.26, 958.4, 962.58, 966.79, 970.97, 975.13, 
    979.24, 983.34, 987.42, 991.46, 995.47, 999.45, 1003.4, 1007.3, 1011.2, 
    1014.9, 1018.7, 1022.5, 1026.4, 1030.2, 1034.1, 1037.9, 1041.7, 1045.4, 
    1049.1, 1052.8, 1056.4, 1060.1, 1063.7, 1067.3, 1070.8, 1074.3, 1077.8, 
    1081.3, 1084.7, 1088.1, 1091.5, 1094.9, 1098.2, 1101.5, 1104.7, 1107.9, 
    1111.1, 1114.2, 1117.4, 1120.5, 1123.6, 1126.7, 1129.8, 1132.9, 1136.1, 
    1139.2, 1142.3, 1145.5, 1148.7, 1151.9, 1155.1, 1158.3, 1161.5, 1164.7, 
    1167.9, 1171.1, 1174.4, 1177.7, 1181, 1184.4, 1187.8, 1191.3, 1194.7, 
    1198.2, 1201.7, 1205.2, 1208.7, 1212.2, 1215.7, 1219.2, 1222.7, 1226.2, 
    1229.7, 1233.1, 1236.6, 1240.1, 1243.5, 1246.9, 1250.4, 1253.9, 1257.4, 
    1260.9, 1264.4, 1268, 1271.5, 1275.1, 1278.6, 1282.2, 1285.6, 1289.1, 
    1292.6, 1296, 1299.4, 1302.7, 1306.1, 1309.4, 1312.6, 1315.8, 1319, 
    1322.1, 1325.3, 1328.4, 1331.5, 1334.6, 1337.8, 1340.9, 1344.1, 1347.3, 
    1350.5, 1353.7, 1357, 1360.2, 1363.5, 1366.8, 1370.1, 1373.4, 1376.7, 
    1380, 1383.3, 1386.6, 1389.9, 1393.1, 1396.4, 1399.6, 1402.8, 1406.1, 
    1409.4, 1412.8, 1416.1, 1419.5, 1422.9, 1426.3, 1429.7, 1433.2, 1436.7, 
    1440.2, 1443.8, 1447.3, 1450.9, 1454.5, 1458.1, 1461.7, 1465.3, 1468.9, 
    1472.5, 1476.1, 1479.7, 1483.3, 1486.9, 1490.5, 1494.1, 1497.8, 1501.4, 
    1505.1, 1508.7, 1512.4, 1516, 1519.7, 1523.3, 1527, 1530.6, 1534.2, 
    1537.9, 1541.5, 1545.1, 1548.7, 1552.2, 1555.8, 1559.4, 1562.9, 1566.5, 
    1570.1, 1573.6, 1577.2, 1580.7, 1584.3, 1587.9, 1591.4, 1595, 1598.6, 
    1602.1, 1605.7, 1609.2, 1612.8, 1616.3, 1619.8, 1623.4, 1626.9, 1630.4, 
    1633.9, 1637.4, 1640.9, 1644.4, 1647.9, 1651.4, 1655, 1658.5, 1662, 
    1665.6, 1669.2, 1672.7, 1676.3, 1679.9, 1683.4, 1687, 1690.5, 1694.1, 
    1697.7, 1701.2, 1704.8, 1708.3, 1711.9, 1715.4, 1718.9, 1722.5, 1726, 
    1729.5, 1733, 1736.6, 1740.1, 1743.6, 1747.2, 1750.7, 1754.3, 1757.8, 
    1761.4, 1764.9, 1768.5, 1772, 1775.5, 1779, 1782.5, 1786, 1789.5, 1793, 
    1796.4, 1799.9, 1803.3, 1806.8, 1810.2, 1813.7, 1817.1, 1820.6, 1824.1, 
    1827.6, 1831.1, 1834.7, 1838.2, 1841.8, 1845.3, 1848.9, 1852.5, 1856, 
    1859.6, 1863.2, 1866.8, 1870.4, 1873.9, 1877.5, 1881.1, 1884.6, 1888.2, 
    1891.8, 1895.3, 1898.9, 1902.5, 1906.1, 1909.6, 1913.2, 1916.8, 1920.4, 
    1924, 1927.7, 1931.3, 1934.9, 1938.5, 1942.2, 1945.8, 1949.4, 1953.1, 
    1956.7, 1960.4, 1964, 1967.6, 1971.2, 1974.8, 1978.4, 1982, 1985.7, 
    1989.3, 1992.9, 1996.5, 2000.1, 2003.8, 2007.4, 2011, 2014.6, 2018.3, 
    2021.9, 2025.5, 2029.1, 2032.8, 2036.4, 2040, 2043.6, 2047.3, 2050.9, 
    2054.5, 2058.1, 2061.7, 2065.3, 2068.9, 2072.5, 2076.1, 2079.7, 2083.3, 
    2086.9, 2090.5, 2094.1, 2097.7, 2101.3, 2104.9, 2108.5, 2112, 2115.6, 
    2119.2, 2122.8, 2126.4, 2130, 2133.6, 2137.2, 2140.8, 2144.4, 2148, 
    2151.6, 2155.2, 2158.9, 2162.5, 2166.2, 2169.9, 2173.5, 2177.2, 2180.9, 
    2184.5, 2188.2, 2191.9, 2195.6, 2199.2, 2202.9, 2206.6, 2210.3, 2213.9, 
    2217.6, 2221.3, 2225, 2228.7, 2232.3, 2236, 2239.7, 2243.4, 2247.1, 
    2250.8, 2254.5, 2258.1, 2261.8, 2265.5, 2269.2, 2272.9, 2276.5, 2280.2, 
    2283.8, 2287.4, 2291, 2294.6, 2298.2, 2301.8, 2305.4, 2308.9, 2312.5, 
    2316.1, 2319.7, 2323.2, 2326.8, 2330.3, 2333.9, 2337.5, 2341, 2344.6, 
    2348.2, 2351.8, 2355.3, 2358.9, 2362.5, 2366.1, 2369.7, 2373.3, 2376.9, 
    2380.5, 2384.1, 2387.7, 2391.2, 2394.8, 2398.3, 2401.9, 2405.4, 2409, 
    2412.5, 2416.1, 2419.6, 2423.1, 2426.7, 2430.2, 2433.7, 2437.2, 2440.8, 
    2444.3, 2447.8, 2451.3, 2454.8, 2458.4, 2461.9, 2465.4, 2469, 2472.5, 
    2476, 2479.5, 2483.1, 2486.6, 2490.1, 2493.6, 2497.1, 2500.6, 2504.1, 
    2507.6, 2511, 2514.5, 2518, 2521.4, 2524.9, 2528.4, 2531.9, 2535.4, 
    2538.9, 2542.4, 2545.9, 2549.4, 2553, 2556.5, 2560.1, 2563.7, 2567.3, 
    2570.9, 2574.5, 2578.2, 2581.8, 2585.4, 2589.1, 2592.8, 2596.4, 2600.1, 
    2603.8, 2607.5, 2611.1, 2614.8, 2618.5, 2622.1, 2625.8, 2629.4, 2633.1, 
    2636.7, 2640.4, 2644, 2647.7, 2651.3, 2655, 2658.6, 2662.3, 2665.9, 
    2669.6, 2673.2, 2676.8, 2680.5, 2684.1, 2687.8, 2691.4, 2695, 2698.6, 
    2702.2, 2705.8, 2709.4, 2713, 2716.5, 2720.1, 2723.7, 2727.2, 2730.8, 
    2734.4, 2737.9, 2741.4, 2745, 2748.5, 2752, 2755.5, 2759.1, 2762.6, 
    2766.1, 2769.6, 2773.1, 2776.7, 2780.2, 2783.7, 2787.2, 2790.8, 2794.3, 
    2797.8, 2801.3, 2804.8, 2808.3, 2811.8, 2815.3, 2818.8, 2822.3, 2825.8, 
    2829.3, 2832.8, 2836.3, 2839.9, 2843.4, 2847, 2850.6, 2854.2, 2857.9, 
    2861.6, 2865.2, 2869, 2872.7, 2876.4, 2880.2, 2884, 2887.8, 2891.6, 
    2895.4, 2899.3, 2903.2, 2907, 2910.9, 2914.9, 2918.8, 2922.8, 2926.8, 
    2930.8, 2934.8, 2938.8, 2942.9, 2947, 2951.1, 2955.2, 2959.3, 2963.5, 
    2967.7, 2971.9, 2976.1, 2980.4, 2984.6, 2988.9, 2993.2, 2997.5, 3001.8, 
    3006.1, 3010.4, 3014.7, 3019, 3023.3, 3027.6, 3031.9, 3036.2, 3040.5, 
    3044.8, 3049.1, 3053.4, 3057.7, 3062, 3066.3, 3070.6, 3074.8, 3079.1, 
    3083.4, 3087.6, 3091.8, 3096.1, 3100.3, 3104.5, 3108.6, 3112.8, 3116.9, 
    3121, 3125.1, 3129.2, 3133.2, 3137.2, 3141.2, 3145.2, 3149.1, 3153, 
    3156.9, 3160.7, 3164.6, 3168.3, 3172.1, 3175.8, 3179.5, 3183.2, 3186.9, 
    3190.6, 3194.2, 3197.9, 3201.5, 3205.1, 3208.7, 3212.3, 3215.8, 3219.4, 
    3223, 3226.5, 3230, 3233.6, 3237.1, 3240.6, 3244.2, 3247.7, 3251.2, 
    3254.7, 3258.3, 3261.8, 3265.3, 3268.9, 3272.4, 3276, 3279.6, 3283.1, 
    3286.7, 3290.2, 3293.8, 3297.4, 3300.9, 3304.5, 3308.1, 3311.6, 3315.2, 
    3318.8, 3322.4, 3325.9, 3329.5, 3333, 3336.6, 3340.2, 3343.7, 3347.2, 
    3350.8, 3354.3, 3357.9, 3361.4, 3364.9, 3368.5, 3372, 3375.6, 3379.1, 
    3382.6, 3386.2, 3389.7, 3393.2, 3396.8, 3400.3, 3403.8, 3407.3, 3410.9, 
    3414.4, 3417.9, 3421.4, 3424.9, 3428.4, 3431.8, 3435.3, 3438.8, 3442.2, 
    3445.7, 3449.1, 3452.6, 3456, 3459.5, 3462.9, 3466.3, 3469.8, 3473.2, 
    3476.6, 3480.1, 3483.5, 3486.9, 3490.4, 3493.8, 3497.2, 3500.6, 3504.1, 
    3507.5, 3510.9, 3514.3, 3517.8, 3521.2, 3524.6, 3528, 3531.4, 3534.8, 
    3538.2, 3541.6, 3545, 3548.4, 3551.8, 3555.2, 3558.6, 3562.1, 3565.5, 
    3568.9, 3572.3, 3575.8, 3579.2, 3582.6, 3586, 3589.5, 3592.9, 3596.3, 
    3599.7, 3603.1, 3606.5, 3609.9, 3613.3, 3616.7, 3620, 3623.4, 3626.8, 
    3630.2, 3633.6, 3637, 3640.4, 3643.8, 3647.3, 3650.7, 3654.1, 3657.5, 
    3660.9, 3664.3, 3667.7, 3671.2, 3674.6, 3678, 3681.4, 3684.8, 3688.3, 
    3691.7, 3695.1, 3698.5, 3701.9, 3705.4, 3708.8, 3712.3, 3715.7, 3719.1, 
    3722.6, 3726, 3729.5, 3733, 3736.4, 3739.9, 3743.4, 3746.9, 3750.4, 
    3753.9, 3757.4, 3760.9, 3764.4, 3767.9, 3771.4, 3774.9, 3778.4, 3781.9, 
    3785.4, 3788.9, 3792.4, 3795.9, 3799.4, 3802.9, 3806.4, 3809.8, 3813.3, 
    3816.8, 3820.3, 3823.8, 3827.2, 3830.7, 3834.2, 3837.7, 3841.1, 3844.6, 
    3848.1, 3851.6, 3855, 3858.5, 3862, 3865.5, 3868.9, 3872.4, 3875.9, 
    3879.3, 3882.8, 3886.2, 3889.7, 3893.1, 3896.6, 3900, 3903.4, 3906.8, 
    3910.2, 3913.7, 3917.1, 3920.5, 3923.9, 3927.3, 3930.7, 3934.2, 3937.6, 
    3941, 3944.4, 3947.9, 3951.3, 3954.7, 3958.2, 3961.6, 3965, 3968.4, 
    3971.9, 3975.3, 3978.7, 3982.1, 3985.5, 3988.9, 3992.3, 3995.8, 3999.2, 
    4002.6, 4006, 4009.4, 4012.9, 4016.3, 4019.7, 4023.1, 4026.6, 4030, 
    4033.4, 4036.9, 4040.3, 4043.7, 4047.2, 4050.6, 4054.1, 4057.5, 4061, 
    4064.4, 4067.9, 4071.3, 4074.8, 4078.3, 4081.7, 4085.2, 4088.7, 4092.2, 
    4095.6, 4099.1, 4102.6, 4106.1, 4109.5, 4113, 4116.5, 4120, 4123.5, 
    4126.9, 4130.4, 4133.9, 4137.4, 4140.9, 4144.3, 4147.8, 4151.3, 4154.7, 
    4158.2, 4161.7, 4165.2, 4168.6, 4172.1, 4175.6, 4179, 4182.5, 4185.9, 
    4189.4, 4192.8, 4196.3, 4199.7, 4203.1, 4206.6, 4210, 4213.4, 4216.8, 
    4220.2, 4223.6, 4227, 4230.4, 4233.8, 4237.2, 4240.6, 4244, 4247.4, 
    4250.8, 4254.2, 4257.6, 4261, 4264.4, 4267.8, 4271.2, 4274.6, 4277.9, 
    4281.3, 4284.7, 4288.1, 4291.5, 4294.9, 4298.2, 4301.6, 4305, 4308.4, 
    4311.8, 4315.2, 4318.5, 4321.9, 4325.3, 4328.7, 4332.1, 4335.5, 4338.9, 
    4342.3, 4345.7, 4349.1, 4352.5, 4355.9, 4359.3, 4362.8, 4366.2, 4369.6, 
    4373, 4376.5, 4379.9, 4383.3, 4386.7, 4390.2, 4393.6, 4397, 4400.4, 
    4403.9, 4407.3, 4410.7, 4414.1, 4417.5, 4421, 4424.4, 4427.8, 4431.3, 
    4434.7, 4438.1, 4441.5, 4445, 4448.4, 4451.8, 4455.3, 4458.7, 4462.1, 
    4465.6, 4469, 4472.5, 4475.9, 4479.4, 4482.8, 4486.2, 4489.7, 4493.1, 
    4496.5, 4500, 4503.4, 4506.8, 4510.2, 4513.7, 4517.1, 4520.5, 4523.9, 
    4527.3, 4530.7, 4534.1, 4537.6, 4541, 4544.4, 4547.8, 4551.2, 4554.6, 
    4558, 4561.4, 4564.8, 4568.2, 4571.6, 4575, 4578.4, 4581.8, 4585.2, 
    4588.6, 4592, 4595.4, 4598.8, 4602.1, 4605.5, 4608.9, 4612.2, 4615.6, 
    4619, 4622.3, 4625.7, 4629, 4632.4, 4635.8, 4639.2, 4642.6, 4646, 4649.3, 
    4652.7, 4656.1, 4659.5, 4662.9, 4666.3, 4669.7, 4673.1, 4676.5, 4679.9, 
    4683.3, 4686.7, 4690.2, 4693.6, 4697, 4700.4, 4703.9, 4707.3, 4710.7, 
    4714.2, 4717.6, 4721, 4724.5, 4727.9, 4731.3, 4734.8, 4738.2, 4741.6, 
    4745.1, 4748.5, 4752, 4755.4, 4758.8, 4762.3, 4765.7, 4769.1, 4772.6, 
    4776, 4779.5, 4782.9, 4786.3, 4789.8, 4793.2, 4796.7, 4800.1, 4803.6, 
    4807, 4810.4, 4813.9, 4817.3, 4820.7, 4824.1, 4827.6, 4831, 4834.4, 
    4837.8, 4841.2, 4844.7, 4848.1, 4851.5, 4855, 4858.4, 4861.8, 4865.3, 
    4868.7, 4872.1, 4875.6, 4879, 4882.4, 4885.8, 4889.3, 4892.7, 4896.1, 
    4899.5, 4902.9, 4906.3, 4909.8, 4913.2, 4916.6, 4920, 4923.4, 4926.8, 
    4930.2, 4933.7, 4937.1, 4940.5, 4943.9, 4947.3, 4950.7, 4954.2, 4957.6, 
    4961, 4964.4, 4967.9, 4971.3, 4974.7, 4978.1, 4981.5, 4985, 4988.4, 
    4991.8, 4995.2, 4998.6, 5002.1, 5005.5, 5008.9, 5012.3, 5015.8, 5019.2, 
    5022.6, 5026.1, 5029.5, 5032.9, 5036.3, 5039.8, 5043.2, 5046.7, 5050.1, 
    5053.5, 5057, 5060.4, 5063.8, 5067.3, 5070.7, 5074.1, 5077.6, 5081, 
    5084.5, 5087.9, 5091.4, 5094.8, 5098.2, 5101.7, 5105.1, 5108.5, 5111.9, 
    5115.3, 5118.8, 5122.2, 5125.6, 5129, 5132.4, 5135.8, 5139.2, 5142.6, 
    5146, 5149.5, 5152.8, 5156.2, 5159.6, 5163, 5166.4, 5169.8, 5173.2, 
    5176.6, 5179.9, 5183.3, 5186.7, 5190, 5193.4, 5196.8, 5200.1, 5203.5, 
    5206.9, 5210.2, 5213.6, 5216.9, 5220.3, 5223.6, 5227, 5230.4, 5233.7, 
    5237.1, 5240.4, 5243.8, 5247.1, 5250.5, 5253.9, 5257.2, 5260.6, 5264, 
    5267.3, 5270.7, 5274, 5277.4, 5280.8, 5284.1, 5287.5, 5290.9, 5294.3, 
    5297.6, 5301, 5304.4, 5307.7, 5311.1, 5314.5, 5317.9, 5321.3, 5324.6, 
    5328, 5331.4, 5334.8, 5338.2, 5341.5, 5344.9, 5348.3, 5351.7, 5355, 
    5358.4, 5361.8, 5365.2, 5368.5, 5371.9, 5375.3, 5378.7, 5382, 5385.4, 
    5388.8, 5392.2, 5395.5, 5398.9, 5402.3, 5405.6, 5409, 5412.4, 5415.7, 
    5419.1, 5422.5, 5425.8, 5429.2, 5432.6, 5435.9, 5439.3, 5442.7, 5446, 
    5449.4, 5452.8, 5456.1, 5459.5, 5462.9, 5466.2, 5469.6, 5473, 5476.4, 
    5479.7, 5483.1, 5486.5, 5489.9, 5493.3, 5496.6, 5500, 5503.4, 5506.8, 
    5510.2, 5513.6, 5517, 5520.3, 5523.7, 5527.1, 5530.5, 5533.9, 5537.3, 
    5540.7, 5544, 5547.4, 5550.8, 5554.2, 5557.6, 5561, 5564.4, 5567.7, 
    5571.1, 5574.5, 5577.9, 5581.2, 5584.6, 5588, 5591.3, 5594.7, 5598, 
    5601.4, 5604.8, 5608.1, 5611.5, 5614.8, 5618.2, 5621.6, 5624.9, 5628.3, 
    5631.6, 5635, 5638.4, 5641.7, 5645.1, 5648.5, 5651.8, 5655.2, 5658.5, 
    5661.9, 5665.2, 5668.6, 5671.9, 5675.3, 5678.6, 5682, 5685.3, 5688.6, 
    5692, 5695.3, 5698.7, 5702.1, 5705.4, 5708.8, 5712.1, 5715.5, 5718.8, 
    5722.2, 5725.6, 5728.9, 5732.3, 5735.6, 5739, 5742.3, 5745.7, 5749, 
    5752.4, 5755.7, 5759.1, 5762.4, 5765.8, 5769.1, 5772.5, 5775.8, 5779.2, 
    5782.5, 5785.9, 5789.2, 5792.6, 5795.9, 5799.3, 5802.6, 5806, 5809.3, 
    5812.7, 5816, 5819.4, 5822.8, 5826.1, 5829.5, 5832.8, 5836.2, 5839.5, 
    5842.9, 5846.2, 5849.6, 5853, 5856.3, 5859.7, 5863, 5866.3, 5869.7, 5873, 
    5876.4, 5879.7, 5883.1, 5886.5, 5889.8, 5893.2, 5896.5, 5899.9, 5903.2, 
    5906.6, 5909.9, 5913.3, 5916.6, 5920, 5923.4, 5926.7, 5930.1, 5933.4, 
    5936.8, 5940.2, 5943.5, 5946.9, 5950.3, 5953.7, 5957, 5960.4, 5963.8, 
    5967.2, 5970.6, 5973.9, 5977.3, 5980.7, 5984.1, 5987.5, 5990.9, 5994.3, 
    5997.6, 6001, 6004.4, 6007.8, 6011.2, 6014.5, 6017.9, 6021.3, 6024.7, 
    6028.1, 6031.5, 6034.8, 6038.2, 6041.6, 6045, 6048.4, 6051.8, 6055.2, 
    6058.6, 6062, 6065.3, 6068.7, 6072.1, 6075.5, 6078.9, 6082.2, 6085.6, 
    6089, 6092.4, 6095.7, 6099.1, 6102.5, 6105.8, 6109.2, 6112.5, 6115.9, 
    6119.2, 6122.6, 6126, 6129.3, 6132.7, 6136.1, 6139.4, 6142.8, 6146.2, 
    6149.5, 6152.9, 6156.2, 6159.6, 6162.9, 6166.3, 6169.6, 6173, 6176.3, 
    6179.6, 6183, 6186.3, 6189.6, 6193, 6196.3, 6199.6, 6203, 6206.3, 6209.6, 
    6213, 6216.3, 6219.7, 6223, 6226.4, 6229.7, 6233, 6236.4, 6239.7, 6243.1, 
    6246.4, 6249.8, 6253.1, 6256.5, 6259.8, 6263.1, 6266.5, 6269.8, 6273.1, 
    6276.5, 6279.8, 6283.2, 6286.5, 6289.9, 6293.2, 6296.5, 6299.9, 6303.2, 
    6306.6, 6310, 6313.3, 6316.7, 6320, 6323.4, 6326.7, 6330.1, 6333.5, 
    6336.8, 6340.2, 6343.5, 6346.9, 6350.2, 6353.6, 6356.9, 6360.3, 6363.6, 
    6367, 6370.3, 6373.7, 6377.1, 6380.4, 6383.8, 6387.1, 6390.5, 6393.9, 
    6397.3, 6400.6, 6404, 6407.4, 6410.7, 6414.1, 6417.5, 6420.8, 6424.2, 
    6427.6, 6431, 6434.3, 6437.7, 6441.1, 6444.5, 6447.9, 6451.2, 6454.6, 
    6458, 6461.4, 6464.8, 6468.1, 6471.5, 6474.9, 6478.3, 6481.7, 6485, 
    6488.4, 6491.8, 6495.2, 6498.6, 6501.9, 6505.3, 6508.7, 6512.1, 6515.5, 
    6518.8, 6522.2, 6525.6, 6529, 6532.3, 6535.7, 6539.1, 6542.5, 6545.8, 
    6549.2, 6552.5, 6555.9, 6559.2, 6562.6, 6565.9, 6569.3, 6572.6, 6576, 
    6579.3, 6582.6, 6586, 6589.3, 6592.6, 6596, 6599.3, 6602.6, 6605.9, 
    6609.3, 6612.6, 6615.9, 6619.2, 6622.5, 6625.8, 6629.2, 6632.5, 6635.8, 
    6639.1, 6642.4, 6645.7, 6649, 6652.2, 6655.5, 6658.8, 6662.1, 6665.4, 
    6668.6, 6671.9, 6675.2, 6678.5, 6681.8, 6685.1, 6688.3, 6691.6, 6694.9, 
    6698.2, 6701.5, 6704.8, 6708, 6711.3, 6714.6, 6717.9, 6721.2, 6724.5, 
    6727.8, 6731.1, 6734.3, 6737.6, 6740.9, 6744.2, 6747.5, 6750.8, 6754.1, 
    6757.4, 6760.7, 6764, 6767.3, 6770.6, 6773.9, 6777.2, 6780.5, 6783.8, 
    6787.1, 6790.5, 6793.8, 6797.1, 6800.4, 6803.7, 6807.1, 6810.4, 6813.7, 
    6817, 6820.3, 6823.7, 6827, 6830.3, 6833.6, 6836.9, 6840.3, 6843.6, 
    6846.9, 6850.2, 6853.6, 6856.9, 6860.2, 6863.5, 6866.9, 6870.2, 6873.5, 
    6876.9, 6880.2, 6883.5, 6886.9, 6890.2, 6893.6, 6896.9, 6900.2, 6903.6, 
    6906.9, 6910.3, 6913.6, 6916.9, 6920.3, 6923.6, 6926.9, 6930.3, 6933.6, 
    6937, 6940.3, 6943.7, 6947, 6950.4, 6953.7, 6957.1, 6960.4, 6963.8, 
    6967.1, 6970.5, 6973.8, 6977.2, 6980.5, 6983.9, 6987.2, 6990.6, 6993.9, 
    6997.3, 7000.6, 7004, 7007.3, 7010.6, 7014, 7017.3, 7020.7, 7024, 7027.4, 
    7030.7, 7034.1, 7037.4, 7040.8, 7044.1, 7047.5, 7050.9, 7054.2, 7057.6, 
    7060.9, 7064.3, 7067.6, 7071, 7074.3, 7077.7, 7081, 7084.3, 7087.7, 7091, 
    7094.3, 7097.7, 7101, 7104.3, 7107.7, 7111, 7114.3, 7117.7, 7121, 7124.4, 
    7127.7, 7131, 7134.4, 7137.7, 7141.1, 7144.4, 7147.7, 7151.1, 7154.4, 
    7157.7, 7161.1, 7164.4, 7167.7, 7171.1, 7174.4, 7177.7, 7181.1, 7184.4, 
    7187.7, 7191, 7194.3, 7197.7, 7201, 7204.3, 7207.7, 7211, 7214.3, 7217.6, 
    7221, 7224.3, 7227.7, 7231, 7234.4, 7237.7, 7241, 7244.4, 7247.7, 7251.1, 
    7254.4, 7257.8, 7261.1, 7264.4, 7267.8, 7271.1, 7274.4, 7277.8, 7281.1, 
    7284.4, 7287.8, 7291.1, 7294.4, 7297.7, 7301.1, 7304.4, 7307.7, 7311.1, 
    7314.4, 7317.8, 7321.1, 7324.4, 7327.8, 7331.1, 7334.4, 7337.8, 7341.1, 
    7344.4, 7347.8, 7351.1, 7354.4, 7357.7, 7361.1, 7364.4, 7367.7, 7371, 
    7374.3, 7377.7, 7381, 7384.3, 7387.6, 7390.9, 7394.2, 7397.5, 7400.9, 
    7404.2, 7407.5, 7410.8, 7414.1, 7417.4, 7420.8, 7424.1, 7427.4, 7430.7, 
    7434, 7437.4, 7440.7, 7444, 7447.3, 7450.6, 7453.9, 7457.2, 7460.5, 
    7463.8, 7467.1, 7470.4, 7473.8, 7477.1, 7480.4, 7483.7, 7487, 7490.3, 
    7493.6, 7497, 7500.3, 7503.6, 7506.9, 7510.2, 7513.5, 7516.8, 7520.1, 
    7523.4, 7526.7, 7530, 7533.3, 7536.6, 7539.9, 7543.2, 7546.5, 7549.8, 
    7553.1, 7556.5, 7559.8, 7563.1, 7566.4, 7569.7, 7573, 7576.4, 7579.7, 
    7583, 7586.3, 7589.6, 7593, 7596.3, 7599.6, 7602.9, 7606.3, 7609.6, 
    7612.9, 7616.2, 7619.5, 7622.8, 7626.2, 7629.5, 7632.8, 7636.1, 7639.4, 
    7642.8, 7646.1, 7649.4, 7652.7, 7656, 7659.3, 7662.7, 7666, 7669.3, 
    7672.6, 7675.9, 7679.3, 7682.6, 7685.9, 7689.2, 7692.5, 7695.9, 7699.2, 
    7702.5, 7705.8, 7709.2, 7712.5, 7715.8, 7719.1, 7722.4, 7725.7, 7729, 
    7732.3, 7735.6, 7738.9, 7742.2, 7745.5, 7748.8, 7752.1, 7755.4, 7758.7, 
    7762, 7765.3, 7768.6, 7771.9, 7775.2, 7778.5, 7781.9, 7785.2, 7788.5, 
    7791.8, 7795.1, 7798.4, 7801.7, 7805, 7808.3, 7811.6, 7814.9, 7818.2, 
    7821.5, 7824.8, 7828.1, 7831.4, 7834.6, 7837.9, 7841.2, 7844.5, 7847.8, 
    7851.1, 7854.4, 7857.7, 7861, 7864.2, 7867.5, 7870.8, 7874.1, 7877.4, 
    7880.7, 7884, 7887.3, 7890.6, 7893.9, 7897.2, 7900.5, 7903.8, 7907, 
    7910.3, 7913.6, 7916.9, 7920.2, 7923.4, 7926.7, 7930, 7933.2, 7936.5, 
    7939.8, 7943.1, 7946.4, 7949.6, 7952.9, 7956.2, 7959.5, 7962.8, 7966, 
    7969.3, 7972.6, 7975.9, 7979.2, 7982.4, 7985.7, 7989, 7992.3, 7995.6, 
    7998.8, 8002.1, 8005.4, 8008.7, 8012, 8015.2, 8018.5, 8021.8, 8025.1, 
    8028.4, 8031.7, 8035, 8038.3, 8041.6, 8044.9, 8048.3, 8051.6, 8054.9, 
    8058.2, 8061.5, 8064.8, 8068.1, 8071.4, 8074.7, 8078, 8081.2, 8084.5, 
    8087.8, 8091.1, 8094.4, 8097.7, 8101, 8104.3, 8107.6, 8110.9, 8114.1, 
    8117.4, 8120.7, 8124, 8127.3, 8130.6, 8133.8, 8137.1, 8140.4, 8143.7, 
    8147, 8150.2, 8153.5, 8156.8, 8160, 8163.3, 8166.6, 8169.8, 8173.1, 
    8176.4, 8179.6, 8182.9, 8186.2, 8189.4, 8192.7, 8195.9, 8199.2, 8202.5, 
    8205.7, 8209, 8212.3, 8215.5, 8218.8, 8222.1, 8225.4, 8228.6, 8231.9, 
    8235.2, 8238.5, 8241.7, 8245, 8248.3, 8251.6, 8254.9, 8258.2, 8261.5, 
    8264.7, 8268, 8271.3, 8274.6, 8277.9, 8281.2, 8284.4, 8287.7, 8291, 
    8294.3, 8297.6, 8300.9, 8304.2, 8307.5, 8310.8, 8314.1, 8317.4, 8320.7, 
    8324, 8327.3, 8330.6, 8333.9, 8337.2, 8340.5, 8343.8, 8347.1, 8350.4, 
    8353.7, 8357, 8360.3, 8363.6, 8366.9, 8370.2, 8373.5, 8376.8, 8380.1, 
    8383.4, 8386.7, 8390, 8393.3, 8396.6, 8399.9, 8403.1, 8406.4, 8409.7, 
    8413, 8416.3, 8419.5, 8422.8, 8426.1, 8429.4, 8432.7, 8436, 8439.3, 
    8442.5, 8445.8, 8449.1, 8452.4, 8455.7, 8459, 8462.2, 8465.5, 8468.8, 
    8472.1, 8475.4, 8478.7, 8481.9, 8485.2, 8488.5, 8491.8, 8495, 8498.3, 
    8501.6, 8504.8, 8508.1, 8511.4, 8514.7, 8517.9, 8521.2, 8524.5, 8527.8, 
    8531.1, 8534.3, 8537.6, 8540.9, 8544.2, 8547.4, 8550.7, 8554, 8557.2, 
    8560.5, 8563.8, 8567, 8570.3, 8573.6, 8576.8, 8580.1, 8583.4, 8586.7, 
    8589.9, 8593.2, 8596.5, 8599.7, 8603, 8606.3, 8609.5, 8612.8, 8616.1, 
    8619.3, 8622.6, 8625.9, 8629.2, 8632.5, 8635.8, 8639, 8642.3, 8645.6, 
    8648.9, 8652.2, 8655.5, 8658.8, 8662.1, 8665.4, 8668.7, 8671.9, 8675.2, 
    8678.5, 8681.8, 8685.1, 8688.4, 8691.7, 8695, 8698.3, 8701.6, 8704.9, 
    8708.2, 8711.5, 8714.8, 8718.1, 8721.4, 8724.7, 8728, 8731.3, 8734.6, 
    8737.9, 8741.2, 8744.5, 8747.8, 8751.1, 8754.4, 8757.7, 8761, 8764.3, 
    8767.6, 8770.9, 8774.2, 8777.4, 8780.7, 8784, 8787.3, 8790.6, 8793.9, 
    8797.2, 8800.5, 8803.8, 8807.1, 8810.4, 8813.7, 8817, 8820.3, 8823.6, 
    8826.9, 8830.1, 8833.4, 8836.7, 8840, 8843.3, 8846.5, 8849.8, 8853, 
    8856.3, 8859.6, 8862.8, 8866.1, 8869.3, 8872.6, 8875.9, 8879.1, 8882.4, 
    8885.6, 8888.9, 8892.2, 8895.4, 8898.7, 8902, 8905.2, 8908.5, 8911.7, 
    8915, 8918.3, 8921.5, 8924.8, 8928, 8931.2, 8934.5, 8937.7, 8941, 8944.2, 
    8947.5, 8950.7, 8954, 8957.2, 8960.5, 8963.7, 8967, 8970.2, 8973.5, 
    8976.8, 8980, 8983.3, 8986.5, 8989.8, 8993, 8996.3, 8999.5, 9002.8, 9006, 
    9009.2, 9012.5, 9015.7, 9019, 9022.2, 9025.5, 9028.7, 9031.9, 9035.2, 
    9038.4, 9041.7, 9044.9, 9048.2, 9051.4, 9054.7, 9057.9, 9061.2, 9064.4, 
    9067.7, 9070.9, 9074.1, 9077.4, 9080.6, 9083.9, 9087.1, 9090.4, 9093.6, 
    9096.9, 9100.1, 9103.4, 9106.6, 9109.9, 9113.1, 9116.4, 9119.6, 9122.9, 
    9126.1, 9129.4, 9132.6, 9135.9, 9139.1, 9142.4, 9145.7, 9148.9, 9152.2, 
    9155.4, 9158.7, 9162, 9165.2, 9168.5, 9171.7, 9175, 9178.2, 9181.5, 
    9184.8, 9188, 9191.3, 9194.6, 9197.8, 9201.1, 9204.3, 9207.6, 9210.9, 
    9214.1, 9217.4, 9220.6, 9223.9, 9227.1, 9230.4, 9233.7, 9236.9, 9240.2, 
    9243.5, 9246.7, 9250, 9253.3, 9256.6, 9259.8, 9263.1, 9266.4, 9269.6, 
    9272.9, 9276.2, 9279.5, 9282.7, 9286, 9289.3, 9292.6, 9295.9, 9299.1, 
    9302.4, 9305.7, 9309, 9312.2, 9315.5, 9318.8, 9322.1, 9325.3, 9328.6, 
    9331.9, 9335.1, 9338.4, 9341.7, 9344.9, 9348.2, 9351.5, 9354.7, 9358, 
    9361.3, 9364.5, 9367.8, 9371.1, 9374.3, 9377.6, 9380.8, 9384.1, 9387.4, 
    9390.6, 9393.9, 9397.1, 9400.4, 9403.7, 9406.9, 9410.2, 9413.4, 9416.7, 
    9420, 9423.2, 9426.5, 9429.7, 9433, 9436.3, 9439.5, 9442.8, 9446.1, 
    9449.3, 9452.6, 9455.9, 9459.1, 9462.4, 9465.7, 9469, 9472.2, 9475.5, 
    9478.8, 9482, 9485.3, 9488.6, 9491.8, 9495.1, 9498.4, 9501.6, 9504.9, 
    9508.2, 9511.4, 9514.7, 9518, 9521.3, 9524.5, 9527.8, 9531.1, 9534.3, 
    9537.6, 9540.9, 9544.1, 9547.4, 9550.7, 9553.9, 9557.2, 9560.5, 9563.8, 
    9567, 9570.3, 9573.6, 9576.8, 9580.1, 9583.4, 9586.6, 9589.9, 9593.2, 
    9596.5, 9599.7, 9603, 9606.3, 9609.6, 9612.8, 9616.1, 9619.4, 9622.7, 
    9625.9, 9629.2, 9632.5, 9635.8, 9639, 9642.3, 9645.6, 9648.8, 9652.1, 
    9655.4, 9658.6, 9661.9, 9665.1, 9668.4, 9671.6, 9674.9, 9678.1, 9681.4, 
    9684.6, 9687.9, 9691.2, 9694.4, 9697.7, 9700.9, 9704.2, 9707.5, 9710.7, 
    9714, 9717.2, 9720.5, 9723.7, 9727, 9730.3, 9733.5, 9736.8, 9740, 9743.2, 
    9746.5, 9749.7, 9753, 9756.2, 9759.5, 9762.7, 9766, 9769.2, 9772.4, 
    9775.7, 9778.9, 9782.2, 9785.4, 9788.7, 9792, 9795.2, 9798.5, 9801.7, 
    9805, 9808.2, 9811.5, 9814.7, 9817.9, 9821.2, 9824.4, 9827.6, 9830.9, 
    9834.1, 9837.4, 9840.6, 9843.9, 9847.1, 9850.3, 9853.6, 9856.8, 9860.1, 
    9863.3, 9866.6, 9869.8, 9873, 9876.3, 9879.5, 9882.7, 9886, 9889.2, 
    9892.5, 9895.7, 9899, 9902.2, 9905.5, 9908.7, 9912, 9915.2, 9918.5, 
    9921.7, 9925, 9928.2, 9931.5, 9934.7, 9938, 9941.2, 9944.5, 9947.7, 
    9950.9, 9954.2, 9957.4, 9960.7, 9963.9, 9967.2, 9970.4, 9973.6, 9976.9, 
    9980.1, 9983.4, 9986.6, 9989.9, 9993.1, 9996.4, 9999.6, 10003, 10006, 
    10009, 10013, 10016, 10019, 10022, 10026, 10029, 10032, 10035, 10039, 
    10042, 10045, 10048, 10052, 10055, 10058, 10061, 10065, 10068, 10071, 
    10074, 10078, 10081, 10084, 10087, 10091, 10094, 10097, 10100, 10104, 
    10107, 10110, 10113, 10116, 10120, 10123, 10126, 10129, 10133, 10136, 
    10139, 10142, 10146, 10149, 10152, 10155, 10159, 10162, 10165, 10168, 
    10172, 10175, 10178, 10181, 10185, 10188, 10191, 10194, 10198, 10201, 
    10204, 10207, 10210, 10214, 10217, 10220, 10223, 10227, 10230, 10233, 
    10236, 10240, 10243, 10246, 10249, 10253, 10256, 10259, 10262, 10266, 
    10269, 10272, 10275, 10279, 10282, 10285, 10288, 10291, 10295, 10298, 
    10301, 10304, 10308, 10311, 10314, 10317, 10320, 10324, 10327, 10330, 
    10333, 10336, 10340, 10343, 10346, 10349, 10353, 10356, 10359, 10362, 
    10365, 10369, 10372, 10375, 10378, 10382, 10385, 10388, 10391, 10395, 
    10398, 10401, 10404, 10408, 10411, 10414, 10417, 10421, 10424, 10427, 
    10430, 10433, 10437, 10440, 10443, 10446, 10450, 10453, 10456, 10460, 
    10463, 10466, 10469, 10473, 10476, 10479, 10482, 10486, 10489, 10492, 
    10495, 10499, 10502, 10505, 10509, 10512, 10515, 10518, 10522, 10525, 
    10528, 10531, 10535, 10538, 10541, 10545, 10548, 10551, 10554, 10558, 
    10561, 10564, 10568, 10571, 10574, 10577, 10581, 10584, 10587, 10591, 
    10594, 10597, 10600, 10604, 10607, 10610, 10614, 10617, 10620, 10623, 
    10627, 10630, 10633, 10637, 10640, 10643, 10647, 10650, 10653, 10656, 
    10660, 10663, 10666, 10670, 10673, 10676, 10679, 10683, 10686, 10689, 
    10693, 10696, 10699, 10702, 10706, 10709, 10712, 10716, 10719, 10722, 
    10726, 10729, 10732, 10736, 10739, 10742, 10745, 10749, 10752, 10755, 
    10759, 10762, 10765, 10769, 10772, 10775, 10779, 10782, 10785, 10788, 
    10792, 10795, 10798, 10802, 10805, 10808, 10812, 10815, 10818, 10822, 
    10825, 10828, 10832, 10835, 10838, 10842, 10845, 10848, 10852, 10855, 
    10858, 10862, 10865, 10868, 10872, 10875, 10878, 10882, 10885, 10888, 
    10891, 10895, 10898, 10901, 10905, 10908, 10911, 10915, 10918, 10921, 
    10925, 10928, 10931, 10935, 10938, 10941, 10945, 10948, 10952, 10955, 
    10958, 10962, 10965, 10968, 10972, 10975, 10978, 10982, 10985, 10988, 
    10991, 10995, 10998, 11001, 11005, 11008, 11011, 11015, 11018, 11021, 
    11025, 11028, 11031, 11034, 11038, 11041, 11044, 11047, 11051, 11054, 
    11057, 11060, 11064, 11067, 11070, 11073, 11077, 11080, 11083, 11086, 
    11089, 11093, 11096, 11099, 11102, 11105, 11109, 11112, 11115, 11118, 
    11122, 11125, 11128, 11131, 11134, 11138, 11141, 11144, 11147, 11151, 
    11154, 11157, 11160, 11164, 11167, 11170, 11173, 11177, 11180, 11183, 
    11186, 11189, 11193, 11196, 11199, 11202, 11206, 11209, 11212, 11215, 
    11218, 11222, 11225, 11228, 11231, 11235, 11238, 11241, 11244, 11247, 
    11251, 11254, 11257, 11260, 11263, 11267, 11270, 11273, 11276, 11280, 
    11283, 11286, 11289, 11292, 11296, 11299, 11302, 11305, 11308, 11312, 
    11315, 11318, 11321, 11325, 11328, 11331, 11334, 11338, 11341, 11344, 
    11347, 11351, 11354, 11357, 11360, 11364, 11367, 11370, 11374, 11377, 
    11380, 11383, 11387, 11390, 11393, 11397, 11400, 11403, 11406, 11410, 
    11413, 11416, 11420, 11423, 11426, 11429, 11433, 11436, 11439, 11443, 
    11446, 11449, 11452, 11456, 11459, 11462, 11466, 11469, 11472, 11475, 
    11479, 11482, 11485, 11488, 11492, 11495, 11498, 11502, 11505, 11508, 
    11511, 11515, 11518, 11521, 11524, 11528, 11531, 11534, 11538, 11541, 
    11544, 11547, 11551, 11554, 11557, 11561, 11564, 11567, 11570, 11574, 
    11577, 11580, 11584, 11587, 11590, 11594, 11597, 11600, 11603, 11607, 
    11610, 11613, 11616, 11620, 11623, 11626, 11630, 11633, 11636, 11639, 
    11643, 11646, 11649, 11653, 11656, 11659, 11662, 11666, 11669, 11672, 
    11675, 11679, 11682, 11685, 11688, 11691, 11695, 11698, 11701, 11704, 
    11708, 11711, 11714, 11718, 11721, 11724, 11727, 11731, 11734, 11737, 
    11741, 11744, 11747, 11750, 11754, 11757, 11760, 11764, 11767, 11770, 
    11773, 11777, 11780, 11783, 11787, 11790, 11793, 11796, 11800, 11803, 
    11806, 11810, 11813, 11816, 11819, 11823, 11826, 11829, 11833, 11836, 
    11839, 11842, 11846, 11849, 11852, 11855, 11859, 11862, 11865, 11869, 
    11872, 11875, 11878, 11882, 11885, 11888, 11891, 11895, 11898, 11901, 
    11905, 11908, 11911, 11914, 11918, 11921, 11924, 11928, 11931, 11934, 
    11937, 11941, 11944, 11947, 11951, 11954, 11957, 11960, 11964, 11967, 
    11970, 11973, 11977, 11980, 11983, 11987, 11990, 11993, 11996, 12000, 
    12003, 12006, 12009, 12013, 12016, 12019, 12022, 12026, 12029, 12032, 
    12035, 12039, 12042, 12045, 12048, 12052, 12055, 12058, 12061, 12065, 
    12068, 12071, 12074, 12078, 12081, 12084, 12087, 12091, 12094, 12097, 
    12100, 12104, 12107, 12110, 12113, 12117, 12120, 12123, 12126, 12130, 
    12133, 12136, 12139, 12142, 12146, 12149, 12152, 12155, 12159, 12162, 
    12165, 12168, 12171, 12175, 12178, 12181, 12184, 12187, 12191, 12194, 
    12197, 12200, 12203, 12207, 12210, 12213, 12216, 12219, 12223, 12226, 
    12229, 12232, 12236, 12239, 12242, 12245, 12249, 12252, 12255, 12258, 
    12261, 12265, 12268, 12271, 12274, 12278, 12281, 12284, 12287, 12291, 
    12294, 12297, 12300, 12304, 12307, 12310, 12313, 12317, 12320, 12323, 
    12326, 12330, 12333, 12336, 12339, 12343, 12346, 12349, 12352, 12355, 
    12359, 12362, 12365, 12368, 12372, 12375, 12378, 12381, 12385, 12388, 
    12391, 12394, 12398, 12401, 12404, 12407, 12411, 12414, 12417, 12420, 
    12424, 12427, 12430, 12433, 12437, 12440, 12443, 12446, 12449, 12453, 
    12456, 12459, 12462, 12466, 12469, 12472, 12475, 12479, 12482, 12485, 
    12488, 12492, 12495, 12498, 12501, 12504, 12508, 12511, 12514, 12517, 
    12520, 12524, 12527, 12530, 12533, 12536, 12540, 12543, 12546, 12549, 
    12553, 12556, 12559, 12562, 12565, 12569, 12572, 12575, 12578, 12581, 
    12585, 12588, 12591, 12594, 12597, 12601, 12604, 12607, 12610, 12613, 
    12617, 12620, 12623, 12626, 12630, 12633, 12636, 12639, 12642, 12646, 
    12649, 12652, 12655, 12659, 12662, 12665, 12668, 12671, 12675, 12678, 
    12681, 12684, 12688, 12691, 12694, 12697, 12700, 12704, 12707, 12710, 
    12713, 12717, 12720, 12723, 12726, 12729, 12733, 12736, 12739, 12742, 
    12746, 12749, 12752, 12755, 12758, 12762, 12765, 12768, 12771, 12774, 
    12778, 12781, 12784, 12787, 12790, 12794, 12797, 12800, 12803, 12806, 
    12810, 12813, 12816, 12819, 12822, 12826, 12829, 12832, 12835, 12838, 
    12842, 12845, 12848, 12851, 12854, 12857, 12861, 12864, 12867, 12870, 
    12873, 12877, 12880, 12883, 12886, 12889, 12893, 12896, 12899, 12902, 
    12913, 12923, 12934, 12944, 12954, 12963, 12973, 12983, 12992, 13002, 
    13011, 13021, 13031, 13041, 13051, 13061, 13072, 13083, 13094, 13105, 
    13117, 13129, 13141, 13154, 13166, 13179, 13192, 13205, 13218, 13232, 
    13245, 13258, 13271, 13284, 13297, 13310, 13322, 13335, 13347, 13359, 
    13371, 13383, 13395, 13406, 13418, 13429, 13441, 13452, 13464, 13476, 
    13487, 13499, 13511, 13522, 13534, 13546, 13559, 13571, 13583, 13596, 
    13608, 13621, 13634, 13646, 13659, 13672, 13685, 13698, 13710, 13723, 
    13736, 13748, 13761, 13773, 13786, 13798, 13811, 13823, 13835, 13847, 
    13859, 13872, 13884, 13896, 13909, 13921, 13933, 13946, 13959, 13971, 
    13984, 13997, 14010, 14023, 14036, 14050, 14063, 14076, 14090, 14103, 
    14117, 14130, 14144, 14157, 14171, 14185, 14198, 14212, 14226, 14239, 
    14253, 14267, 14280, 14294, 14307, 14321, 14334, 14348, 14362, 14375, 
    14388, 14402, 14415, 14428, 14442, 14455, 14468, 14481, 14495, 14508, 
    14521, 14534, 14547, 14560, 14573, 14586, 14599, 14612, 14625, 14639, 
    14652, 14665, 14678, 14692, 14705, 14719, 14733, 14747, 14761, 14775, 
    14789, 14804, 14818, 14833, 14848, 14863, 14878, 14893, 14908, 14924, 
    14939, 14955, 14971, 14986, 15002, 15018, 15034, 15049, 15065, 15081, 
    15097, 15113, 15129, 15144, 15160, 15176, 15192, 15208, 15223, 15239, 
    15255, 15271, 15286, 15302, 15318, 15333, 15349, 15365, 15380, 15396, 
    15412, 15427, 15443, 15459, 15475, 15490, 15506, 15522, 15538, 15553, 
    15569, 15585, 15601, 15618, 15634, 15650, 15667, 15684, 15701, 15718, 
    15736, 15753, 15772, 15790, 15808, 15827, 15846, 15866, 15885, 15905, 
    15925, 15945, 15966, 15986, 16007, 16028, 16048, 16069, 16090, 16111, 
    16132, 16152, 16173, 16194, 16215, 16235, 16256, 16277, 16297, 16318, 
    16338, 16359, 16379, 16400, 16420, 16440, 16460, 16481, 16501, 16521, 
    16540, 16560, 16580, 16599, 16618, 16637, 16656, 16675, 16693, 16711, 
    16729, 16746, 16764, 16781, 16798, 16814, 16831, 16847, 16863, 16878, 
    16894, 16909, 16925, 16940, 16955, 16970, 16985, 17000, 17015, 17030, 
    17046, 17061, 17076, 17092, 17107, 17122, 17138, 17153, 17169, 17185, 
    17200, 17216, 17232, 17247, 17263, 17279, 17295, 17310, 17326, 17342, 
    17358, 17375, 17391, 17408, 17424, 17441, 17458, 17476, 17493, 17511, 
    17529, 17547, 17566, 17585, 17604, 17623, 17642, 17662, 17682, 17702, 
    17723, 17743, 17764, 17785, 17806, 17828, 17849, 17871, 17893, 17915, 
    17937, 17959, 17982, 18004, 18027, 18049, 18072, 18095, 18118, 18141, 
    18163, 18186, 18209, 18232, 18254, 18277, 18300, 18322, 18345, 18367, 
    18389, 18412, 18434, 18456, 18478, 18499, 18521, 18543, 18564, 18585, 
    18606, 18628, 18648, 18669, 18690, 18711, 18731, 18752, 18772, 18792, 
    18812, 18832, 18852, 18872, 18892, 18912, 18931, 18951, 18971, 18990, 
    19010, 19029, 19049, 19068, 19088, 19107, 19127, 19146, 19166, 19185, 
    19204, 19224, 19243, 19262, 19282, 19301, 19320, 19340, 19359, 19379, 
    19398, 19418, 19438, 19458, 19478, 19498, 19519, 19539, 19560, 19581, 
    19602, 19624, 19645, 19667, 19689, 19711, 19733, 19755, 19777, 19799, 
    19822, 19844, 19866, 19889, 19911, 19933, 19955, 19977, 19999, 20021, 
    20043, 20065, 20087, 20108, 20130, 20152, 20173, 20195, 20217, 20238, 
    20260, 20282, 20304, 20326, 20348, 20370, 20392, 20414, 20436, 20459, 
    20481, 20503, 20526, 20548, 20571, 20593, 20616, 20639, 20662, 20685, 
    20708, 20731, 20754, 20778, 20801, 20825, 20849, 20874, 20898, 20923, 
    20948, 20973, 20998, 21024, 21049, 21075, 21101, 21127, 21153, 21180, 
    21206, 21232, 21259, 21285, 21311, 21337, 21363, 21389, 21415, 21441, 
    21467, 21492, 21517, 21542, 21567, 21592, 21616, 21640, 21664, 21688, 
    21712, 21735, 21758, 21781, 21804, 21827, 21849, 21872, 21894, 21916, 
    21939, 21961, 21984, 22006, 22029, 22052, 22075, 22098, 22121, 22145, 
    22169, 22193, 22218, 22243, 22268, 22294, 22319, 22346, 22372, 22399, 
    22425, 22453, 22480, 22507, 22535, 22563, 22591, 22619, 22647, 22675, 
    22703, 22731, 22759, 22787, 22815, 22843, 22871, 22898, 22926, 22954, 
    22982, 23009, 23037, 23064, 23092, 23120, 23147, 23175, 23202, 23230, 
    23257, 23285, 23312, 23339, 23366, 23394, 23421, 23448, 23474, 23501, 
    23527, 23554, 23580, 23606, 23631, 23657, 23683, 23708, 23733, 23758, 
    23783, 23808, 23833, 23858, 23883, 23908, 23934, 23959, 23984, 24010, 
    24035, 24061, 24087, 24113, 24140, 24166, 24193, 24220, 24247, 24275, 
    24302, 24330, 24358, 24387, 24415, 24444, 24473, 24502, 24532, 24561, 
    24591, 24621, 24651, 24682, 24712, 24743, 24773, 24804, 24835, 24865, 
    24896, 24927, 24957, 24988, 25019, 25049, 25080, 25110, 25141, 25171, 
    25202, 25232, 25262, 25292, 25323, 25353, 25383, 25413, 25443, 25473, 
    25503, 25533, 25562, 25592, 25622, 25651, 25681, 25711, 25740, 25770, 
    25799, 25829, 25858, 25887, 25917, 25946, 25976, 26005, 26035, 26064, 
    26094, 26123, 26153, 26182, 26211, 26240, 26269, 26298, 26326, 26355, 
    26383, 26412, 26440, 26468, 26496, 26525, 26553, 26581, 26610, 26638, 
    26667, 26696, 26725, 26754, 26783, 26813, 26843, 26873, 26903, 26933, 
    26964, 26995, 27026, 27058, 27090, 27122, 27154, 27186, 27219, 27252, 
    27285, 27318, 27351, 27385, 27419, 27452, 27486, 27520, 27554, 27588, 
    27622, 27656, 27689, 27723, 27757, 27790, 27824, 27857, 27890, 27923, 
    27956, 27989, 28022, 28055, 28087, 28120, 28153, 28185, 28217, 28250, 
    28282, 28314, 28346, 28378, 28410, 28442, 28474, 28506, 28539, 28571, 
    28603, 28635, 28667, 28699, 28731, 28763, 28795, 28827, 28859, 28891, 
    28923, 28956, 28988, 29020, 29052, 29084, 29116, 29148, 29180, 29212, 
    29244, 29276, 29308, 29340, 29372, 29404, 29436, 29468, 29499, 29531, 
    29563, 29594, 29626, 29657, 29689, 29720, 29752, 29783, 29814, 29846, 
    29877, 29909, 29940, 29972, 30004, 30036, 30068, 30100, 30132, 30165, 
    30198, 30230, 30263, 30297, 30330, 30364, 30397, 30431, 30465, 30499, 
    30534, 30568, 30603, 30637, 30672, 30706, 30741, 30776, 30810, 30845, 
    30879, 30914, 30949, 30983, 31018, 31052, 31087, 31121, 31155, 31190, 
    31224, 31258, 31292, 31327, 31361, 31395, 31429, 31463, 31497, 31531, 
    31566, 31600, 31634, 31668, 31703, 31737, 31772, 31806, 31841, 31875, 
    31910, 31945, 31980, 32015, 32050, 32085, 32120, 32155, 32191, 32226, 
    32261, 32296, 32331, 32367, 32402, 32437, 32472, 32507, 32543, 32578, 
    32613, 32648, 32683, 32718, 32753, 32789, 32824, 32859, 32894, 32929, 
    32965, 33000, 33036, 33071, 33107, 33142, 33178, 33213, 33249, 33285, 
    33320, 33356, 33392, 33427, 33463, 33499, 33534, 33570, 33606, 33641, 
    33677, 33712, 33748, 33783, 33818, 33854, 33889, 33924, 33959, 33994, 
    34030, 34065, 34100, 34135, 34170, 34205, 34240, 34274, 34309, 34344, 
    34379, 34414, 34449, 34484, 34519, 34554, 34589, 34624, 34659, 34694, 
    34729, 34764, 34799, 34835, 34870, 34905, 34940, 34976, 35011, 35047, 
    35083, 35118, 35154, 35190, 35226, 35262, 35298, 35334, 35370, 35406, 
    35442, 35478, 35514, 35550, 35586, 35622, 35658, 35694, 35730, 35765, 
    35801, 35837, 35872, 35908, 35943, 35979, 36014, 36050, 36086, 36121, 
    36157, 36193, 36229, 36265, 36301, 36337, 36373, 36410, 36446, 36482, 
    36519, 36555, 36592, 36629, 36665, 36702, 36738, 36775, 36812, 36848, 
    36885, 36921, 36957, 36994, 37030, 37066, 37102, 37139, 37175, 37210, 
    37246, 37282, 37318, 37353, 37389, 37424, 37460, 37495, 37531, 37566, 
    37601, 37636, 37672, 37707, 37742, 37777, 37813, 37848, 37884, 37919, 
    37955, 37990, 38026, 38062, 38098, 38134, 38170, 38206, 38242, 38279, 
    38315, 38352, 38388, 38425, 38462, 38499, 38536, 38573, 38611, 38648, 
    38685, 38723, 38760, 38797, 38835, 38872, 38910, 38947, 38984, 39022, 
    39059, 39096, 39133, 39170, 39207, 39244, 39281, 39318, 39355, 39392, 
    39429, 39465, 39502, 39539, 39575, 39612, 39649, 39685, 39722, 39758, 
    39795, 39831, 39868, 39904, 39940, 39977, 40013, 40049, 40086, 40122, 
    40158, 40194, 40231, 40267, 40303, 40339, 40376, 40412, 40448, 40485, 
    40521, 40557, 40594, 40630, 40667, 40703, 40740, 40776, 40813, 40849, 
    40886, 40922, 40959, 40995, 41032, 41068, 41105, 41142, 41178, 41215, 
    41252, 41288, 41325, 41362, 41398, 41435, 41472, 41509, 41546, 41583, 
    41619, 41656, 41693, 41730, 41767, 41804, 41841, 41878, 41915, 41952, 
    41989, 42026, 42062, 42099, 42136, 42173, 42210, 42247, 42284, 42321, 
    42357, 42394, 42431, 42468, 42505, 42542, 42578, 42615, 42652, 42689, 
    42725, 42762, 42799, 42836, 42873, 42909, 42946, 42983, 43020, 43057, 
    43094, 43131, 43168, 43205, 43242, 43279, 43316, 43354, 43391, 43428, 
    43466, 43503, 43540, 43578, 43615, 43652, 43690, 43727, 43765, 43802, 
    43840, 43877, 43914, 43952, 43989, 44027, 44064, 44101, 44139, 44176, 
    44213, 44251, 44288, 44325, 44362, 44399, 44436, 44473, 44511, 44548, 
    44585, 44622, 44659, 44696, 44733, 44770, 44808, 44845, 44882, 44920, 
    44957, 44995, 45033, 45071, 45108, 45146, 45184, 45222, 45260, 45298, 
    45336, 45374, 45412, 45450, 45487, 45525, 45562, 45599, 45636, 45673, 
    45709, 45746, 45782, 45818, 45854, 45890, 45926, 45962, 45997, 46033, 
    46068, 46104, 46140, 46175, 46211, 46246, 46282, 46318, 46354, 46390, 
    46427, 46463, 46500, 46536, 46573, 46611, 46648, 46685, 46723, 46760, 
    46798, 46836, 46874, 46912, 46950, 46988, 47026, 47065, 47103, 47141, 
    47179, 47217, 47255, 47293, 47331, 47369, 47407, 47445, 47482, 47520, 
    47557, 47594, 47631, 47668, 47705, 47741, 47778, 47814, 47851, 47887, 
    47923, 47959, 47996, 48032, 48068, 48104, 48140, 48176, 48212, 48248, 
    48284, 48321, 48357, 48393, 48430, 48466, 48502, 48539, 48575, 48612, 
    48648, 48685, 48721, 48758, 48794, 48831, 48868, 48905, 48941, 48978, 
    49015, 49052, 49089, 49127, 49164, 49201, 49239, 49276, 49314, 49352, 
    49389, 49427, 49465, 49503, 49541, 49579, 49617, 49655, 49693, 49731, 
    49769, 49807, 49845, 49883, 49921, 49958, 49996, 50034, 50071, 50109, 
    50146, 50184, 50221, 50258, 50296, 50333, 50370, 50407, 50445, 50482, 
    50519, 50556, 50594, 50631, 50668, 50705, 50742, 50779, 50817, 50854, 
    50891, 50927, 50964, 51001, 51038, 51075, 51111, 51148, 51184, 51221, 
    51257, 51294, 51330, 51367, 51403, 51440, 51476, 51513, 51549, 51586, 
    51622, 51659, 51696, 51732, 51769, 51805, 51842, 51879, 51915, 51952, 
    51988, 52024, 52061, 52097, 52133, 52170, 52206, 52242, 52278, 52314, 
    52350, 52386, 52422, 52458, 52495, 52531, 52567, 52603, 52639, 52675, 
    52712, 52748, 52784, 52821, 52857, 52894, 52930, 52967, 53003, 53040, 
    53076, 53113, 53149, 53186, 53223, 53259, 53296, 53333, 53370, 53407, 
    53444, 53481, 53518, 53555, 53592, 53629, 53667, 53704, 53741, 53779, 
    53816, 53853, 53890, 53927, 53965, 54002, 54039, 54076, 54113, 54150, 
    54187, 54223, 54260, 54297, 54334, 54371, 54407, 54444, 54481, 54518, 
    54554, 54591, 54628, 54665, 54701, 54738, 54775, 54812, 54849, 54886, 
    54923, 54960, 54996, 55033, 55070, 55107, 55144, 55181, 55218, 55255, 
    55292, 55329, 55366, 55403, 55440, 55477, 55514, 55551, 55587, 55624, 
    55661, 55698, 55735, 55772, 55809, 55846, 55883, 55919, 55956, 55993, 
    56030, 56066, 56103, 56140, 56176, 56213, 56249, 56286, 56323, 56359, 
    56396, 56432, 56469, 56505, 56542, 56579, 56615, 56652, 56689, 56726, 
    56763, 56800, 56837, 56875, 56912, 56950, 56987, 57025, 57062, 57100, 
    57138, 57176, 57214, 57251, 57289, 57327, 57364, 57402, 57440, 57477, 
    57514, 57551, 57589, 57626, 57663, 57699, 57736, 57773, 57809, 57846, 
    57883, 57919, 57956, 57992, 58028, 58065, 58101, 58138, 58174, 58211, 
    58247, 58284, 58320, 58357, 58393, 58430, 58467, 58503, 58540, 58576, 
    58613, 58650, 58686, 58723, 58759, 58796, 58833, 58869, 58906, 58943, 
    58979, 59016, 59053, 59089, 59126, 59163, 59199, 59236, 59273, 59310, 
    59347, 59383, 59420, 59457, 59494, 59531, 59568, 59605, 59643, 59680, 
    59717, 59754, 59791, 59829, 59866, 59903, 59941, 59978 ;

 geop_refrac =
  31.017, 32.515, 33.964, 35.36, 36.725, 38.09, 39.472, 40.889, 42.331, 
    43.799, 45.325, 46.934, 48.636, 50.438, 52.35, 54.39, 56.578, 58.889, 
    61.33, 63.893, 66.584, 69.407, 72.337, 75.365, 78.42, 81.509, 84.638, 
    87.821, 91.059, 94.324, 97.614, 100.92, 104.27, 107.67, 111.12, 114.65, 
    118.24, 121.9, 125.62, 129.38, 133.19, 137.02, 140.9, 144.82, 148.76, 
    152.72, 156.67, 160.61, 164.52, 168.43, 172.33, 176.23, 180.12, 183.99, 
    187.85, 191.68, 195.5, 199.3, 203.07, 206.84, 210.64, 214.45, 218.29, 
    222.17, 226.06, 229.95, 233.82, 237.68, 241.54, 245.4, 249.26, 253.1, 
    256.93, 260.72, 264.48, 268.2, 271.91, 275.6, 279.3, 282.98, 286.65, 
    290.29, 293.9, 297.52, 301.16, 304.83, 308.51, 312.2, 315.91, 319.63, 
    323.35, 327.08, 330.84, 334.61, 338.41, 342.23, 346.05, 349.89, 353.74, 
    357.6, 361.47, 365.34, 369.22, 373.1, 376.98, 380.88, 384.79, 388.7, 
    392.63, 396.55, 400.47, 404.39, 408.32, 412.26, 416.21, 420.16, 424.1, 
    428.05, 431.99, 435.92, 439.83, 443.72, 447.6, 451.47, 455.32, 459.17, 
    463, 466.82, 470.63, 474.44, 478.25, 482.06, 485.86, 489.65, 493.45, 
    497.26, 501.06, 504.88, 508.7, 512.53, 516.36, 520.19, 524.02, 527.85, 
    531.69, 535.53, 539.36, 543.18, 547.02, 550.85, 554.69, 558.53, 562.36, 
    566.18, 570.01, 573.86, 577.72, 581.58, 585.45, 589.35, 593.27, 597.22, 
    601.21, 605.21, 609.24, 613.29, 617.37, 621.46, 625.58, 629.71, 633.88, 
    638.07, 642.29, 646.53, 650.78, 655.05, 659.34, 663.65, 667.99, 672.37, 
    676.78, 681.24, 685.73, 690.28, 694.89, 699.58, 704.36, 709.23, 714.18, 
    719.23, 724.39, 729.67, 735, 740.38, 745.76, 751.14, 756.52, 761.89, 
    767.25, 772.56, 777.83, 783.05, 788.28, 793.51, 798.75, 803.99, 809.24, 
    814.51, 819.79, 825.05, 830.3, 835.55, 840.8, 846.06, 851.3, 856.5, 
    861.61, 866.66, 871.66, 876.63, 881.56, 886.45, 891.28, 896.05, 900.72, 
    905.3, 909.77, 914.12, 918.36, 922.52, 926.61, 930.63, 934.63, 938.63, 
    942.66, 946.7, 950.76, 954.85, 958.99, 963.17, 967.38, 971.57, 975.73, 
    979.84, 983.94, 988.02, 992.07, 996.08, 1000.1, 1004, 1007.9, 1011.8, 
    1015.6, 1019.3, 1023.1, 1027, 1030.8, 1034.7, 1038.5, 1042.3, 1046.1, 
    1049.8, 1053.4, 1057.1, 1060.7, 1064.3, 1067.9, 1071.4, 1075, 1078.5, 
    1081.9, 1085.4, 1088.8, 1092.2, 1095.5, 1098.9, 1102.1, 1105.4, 1108.5, 
    1111.7, 1114.9, 1118, 1121.2, 1124.3, 1127.4, 1130.5, 1133.6, 1136.7, 
    1139.9, 1143, 1146.2, 1149.4, 1152.6, 1155.8, 1159, 1162.2, 1165.4, 
    1168.6, 1171.8, 1175, 1178.4, 1181.7, 1185.1, 1188.5, 1192, 1195.4, 
    1198.9, 1202.4, 1205.9, 1209.4, 1212.9, 1216.4, 1219.9, 1223.4, 1226.9, 
    1230.4, 1233.8, 1237.3, 1240.8, 1244.2, 1247.7, 1251.1, 1254.6, 1258.1, 
    1261.6, 1265.2, 1268.7, 1272.3, 1275.8, 1279.4, 1282.9, 1286.4, 1289.8, 
    1293.3, 1296.7, 1300.1, 1303.5, 1306.8, 1310.1, 1313.4, 1316.6, 1319.7, 
    1322.9, 1326, 1329.1, 1332.2, 1335.4, 1338.5, 1341.7, 1344.8, 1348, 
    1351.2, 1354.5, 1357.7, 1361, 1364.2, 1367.5, 1370.9, 1374.2, 1377.5, 
    1380.8, 1384.1, 1387.4, 1390.6, 1393.9, 1397.1, 1400.3, 1403.6, 1406.9, 
    1410.2, 1413.5, 1416.9, 1420.2, 1423.6, 1427.1, 1430.5, 1434, 1437.5, 
    1441, 1444.5, 1448.1, 1451.7, 1455.3, 1458.9, 1462.5, 1466.1, 1469.7, 
    1473.3, 1476.9, 1480.5, 1484.1, 1487.7, 1491.3, 1494.9, 1498.6, 1502.2, 
    1505.9, 1509.5, 1513.2, 1516.8, 1520.5, 1524.1, 1527.8, 1531.4, 1535, 
    1538.7, 1542.3, 1545.9, 1549.5, 1553, 1556.6, 1560.2, 1563.8, 1567.3, 
    1570.9, 1574.4, 1578, 1581.6, 1585.1, 1588.7, 1592.3, 1595.8, 1599.4, 
    1602.9, 1606.5, 1610, 1613.6, 1617.1, 1620.7, 1624.2, 1627.7, 1631.2, 
    1634.7, 1638.2, 1641.8, 1645.3, 1648.8, 1652.3, 1655.8, 1659.3, 1662.9, 
    1666.4, 1670, 1673.6, 1677.1, 1680.7, 1684.3, 1687.8, 1691.4, 1695, 
    1698.5, 1702.1, 1705.6, 1709.2, 1712.7, 1716.3, 1719.8, 1723.3, 1726.9, 
    1730.4, 1733.9, 1737.4, 1740.9, 1744.5, 1748, 1751.6, 1755.1, 1758.7, 
    1762.2, 1765.8, 1769.3, 1772.8, 1776.4, 1779.9, 1783.4, 1786.9, 1790.4, 
    1793.8, 1797.3, 1800.7, 1804.2, 1807.6, 1811.1, 1814.5, 1818, 1821.5, 
    1825, 1828.5, 1832, 1835.5, 1839.1, 1842.6, 1846.2, 1849.8, 1853.3, 
    1856.9, 1860.5, 1864.1, 1867.7, 1871.2, 1874.8, 1878.4, 1882, 1885.5, 
    1889.1, 1892.6, 1896.2, 1899.8, 1903.4, 1906.9, 1910.5, 1914.1, 1917.7, 
    1921.3, 1924.9, 1928.5, 1932.2, 1935.8, 1939.4, 1943.1, 1946.7, 1950.3, 
    1954, 1957.6, 1961.2, 1964.9, 1968.5, 1972.1, 1975.7, 1979.3, 1982.9, 
    1986.6, 1990.2, 1993.8, 1997.4, 2001, 2004.7, 2008.3, 2011.9, 2015.5, 
    2019.2, 2022.8, 2026.4, 2030.1, 2033.7, 2037.3, 2040.9, 2044.5, 2048.2, 
    2051.8, 2055.4, 2059, 2062.6, 2066.2, 2069.8, 2073.4, 2077, 2080.7, 
    2084.2, 2087.8, 2091.4, 2095, 2098.6, 2102.2, 2105.8, 2109.4, 2113, 
    2116.5, 2120.1, 2123.7, 2127.3, 2130.9, 2134.5, 2138.1, 2141.7, 2145.3, 
    2148.9, 2152.5, 2156.2, 2159.8, 2163.5, 2167.1, 2170.8, 2174.4, 2178.1, 
    2181.8, 2185.4, 2189.1, 2192.8, 2196.5, 2200.2, 2203.8, 2207.5, 2211.2, 
    2214.9, 2218.5, 2222.2, 2225.9, 2229.6, 2233.3, 2236.9, 2240.6, 2244.3, 
    2248, 2251.7, 2255.4, 2259.1, 2262.8, 2266.4, 2270.1, 2273.8, 2277.4, 
    2281.1, 2284.7, 2288.3, 2291.9, 2295.6, 2299.1, 2302.7, 2306.3, 2309.9, 
    2313.5, 2317, 2320.6, 2324.2, 2327.7, 2331.3, 2334.8, 2338.4, 2342, 
    2345.5, 2349.1, 2352.7, 2356.3, 2359.9, 2363.5, 2367, 2370.6, 2374.2, 
    2377.8, 2381.4, 2385, 2388.6, 2392.2, 2395.7, 2399.3, 2402.8, 2406.4, 
    2409.9, 2413.4, 2417, 2420.5, 2424.1, 2427.6, 2431.1, 2434.6, 2438.2, 
    2441.7, 2445.2, 2448.7, 2452.3, 2455.8, 2459.3, 2462.8, 2466.4, 2469.9, 
    2473.4, 2476.9, 2480.5, 2484, 2487.5, 2491, 2494.6, 2498.1, 2501.5, 2505, 
    2508.5, 2512, 2515.4, 2518.9, 2522.4, 2525.8, 2529.3, 2532.8, 2536.3, 
    2539.8, 2543.3, 2546.8, 2550.3, 2553.9, 2557.4, 2561, 2564.6, 2568.2, 
    2571.8, 2575.5, 2579.1, 2582.7, 2586.4, 2590, 2593.7, 2597.4, 2601, 
    2604.7, 2608.4, 2612.1, 2615.7, 2619.4, 2623.1, 2626.7, 2630.3, 2634, 
    2637.6, 2641.3, 2644.9, 2648.6, 2652.2, 2655.9, 2659.6, 2663.2, 2666.8, 
    2670.5, 2674.1, 2677.8, 2681.4, 2685, 2688.7, 2692.3, 2695.9, 2699.5, 
    2703.1, 2706.7, 2710.3, 2713.9, 2717.5, 2721, 2724.6, 2728.2, 2731.7, 
    2735.3, 2738.8, 2742.3, 2745.9, 2749.4, 2752.9, 2756.4, 2760, 2763.5, 
    2767, 2770.5, 2774.1, 2777.6, 2781.1, 2784.6, 2788.1, 2791.7, 2795.2, 
    2798.7, 2802.2, 2805.7, 2809.2, 2812.8, 2816.2, 2819.7, 2823.2, 2826.7, 
    2830.2, 2833.7, 2837.2, 2840.8, 2844.3, 2847.9, 2851.5, 2855.1, 2858.8, 
    2862.5, 2866.2, 2869.9, 2873.6, 2877.3, 2881.1, 2884.9, 2888.7, 2892.5, 
    2896.3, 2900.2, 2904.1, 2907.9, 2911.8, 2915.8, 2919.7, 2923.7, 2927.7, 
    2931.7, 2935.7, 2939.7, 2943.8, 2947.8, 2951.9, 2956.1, 2960.2, 2964.4, 
    2968.6, 2972.8, 2977, 2981.3, 2985.5, 2989.8, 2994.1, 2998.4, 3002.7, 
    3007, 3011.2, 3015.5, 3019.8, 3024.1, 3028.5, 3032.8, 3037.1, 3041.4, 
    3045.7, 3049.9, 3054.2, 3058.5, 3062.8, 3067.1, 3071.4, 3075.7, 3080, 
    3084.2, 3088.5, 3092.7, 3096.9, 3101.1, 3105.3, 3109.5, 3113.6, 3117.8, 
    3121.9, 3126, 3130, 3134.1, 3138.1, 3142.1, 3146, 3150, 3153.9, 3157.7, 
    3161.6, 3165.4, 3169.2, 3172.9, 3176.7, 3180.4, 3184.1, 3187.7, 3191.4, 
    3195.1, 3198.7, 3202.3, 3205.9, 3209.5, 3213.1, 3216.7, 3220.2, 3223.8, 
    3227.3, 3230.9, 3234.4, 3237.9, 3241.5, 3245, 3248.5, 3252, 3255.6, 
    3259.1, 3262.6, 3266.2, 3269.7, 3273.3, 3276.8, 3280.4, 3283.9, 3287.5, 
    3291.1, 3294.6, 3298.2, 3301.8, 3305.3, 3308.9, 3312.5, 3316, 3319.6, 
    3323.2, 3326.7, 3330.3, 3333.9, 3337.4, 3341, 3344.5, 3348, 3351.6, 
    3355.1, 3358.7, 3362.2, 3365.7, 3369.3, 3372.8, 3376.4, 3379.9, 3383.4, 
    3387, 3390.5, 3394, 3397.6, 3401.1, 3404.6, 3408.1, 3411.6, 3415.1, 
    3418.6, 3422.1, 3425.6, 3429.1, 3432.6, 3436.1, 3439.5, 3443, 3446.4, 
    3449.9, 3453.3, 3456.8, 3460.2, 3463.7, 3467.1, 3470.5, 3473.9, 3477.4, 
    3480.8, 3484.2, 3487.7, 3491.1, 3494.5, 3498, 3501.4, 3504.8, 3508.2, 
    3511.7, 3515.1, 3518.5, 3521.9, 3525.3, 3528.7, 3532.1, 3535.5, 3538.9, 
    3542.3, 3545.8, 3549.2, 3552.6, 3556, 3559.4, 3562.8, 3566.2, 3569.6, 
    3573.1, 3576.5, 3579.9, 3583.3, 3586.8, 3590.2, 3593.6, 3597, 3600.4, 
    3603.8, 3607.2, 3610.6, 3614, 3617.4, 3620.8, 3624.2, 3627.5, 3630.9, 
    3634.3, 3637.7, 3641.1, 3644.5, 3648, 3651.4, 3654.8, 3658.2, 3661.6, 
    3665, 3668.4, 3671.8, 3675.3, 3678.7, 3682.1, 3685.5, 3688.9, 3692.4, 
    3695.8, 3699.2, 3702.6, 3706.1, 3709.5, 3712.9, 3716.4, 3719.8, 3723.3, 
    3726.7, 3730.2, 3733.6, 3737.1, 3740.6, 3744.1, 3747.6, 3751, 3754.5, 
    3758, 3761.5, 3765, 3768.5, 3772, 3775.5, 3779, 3782.5, 3786, 3789.5, 
    3793, 3796.5, 3800, 3803.5, 3807, 3810.5, 3814, 3817.4, 3820.9, 3824.4, 
    3827.9, 3831.3, 3834.8, 3838.3, 3841.8, 3845.2, 3848.7, 3852.2, 3855.7, 
    3859.1, 3862.6, 3866.1, 3869.5, 3873, 3876.5, 3879.9, 3883.4, 3886.8, 
    3890.3, 3893.7, 3897.2, 3900.6, 3904, 3907.4, 3910.8, 3914.2, 3917.7, 
    3921.1, 3924.5, 3927.9, 3931.3, 3934.7, 3938.2, 3941.6, 3945, 3948.4, 
    3951.9, 3955.3, 3958.7, 3962.1, 3965.6, 3969, 3972.4, 3975.8, 3979.3, 
    3982.7, 3986.1, 3989.5, 3992.9, 3996.3, 3999.7, 4003.1, 4006.6, 4010, 
    4013.4, 4016.8, 4020.2, 4023.7, 4027.1, 4030.5, 4033.9, 4037.4, 4040.8, 
    4044.3, 4047.7, 4051.1, 4054.6, 4058, 4061.5, 4064.9, 4068.4, 4071.8, 
    4075.3, 4078.8, 4082.2, 4085.7, 4089.2, 4092.7, 4096.1, 4099.6, 4103.1, 
    4106.6, 4110, 4113.5, 4117, 4120.5, 4123.9, 4127.4, 4130.9, 4134.4, 
    4137.9, 4141.3, 4144.8, 4148.3, 4151.7, 4155.2, 4158.7, 4162.2, 4165.6, 
    4169.1, 4172.5, 4176, 4179.5, 4182.9, 4186.4, 4189.8, 4193.3, 4196.7, 
    4200.1, 4203.6, 4207, 4210.4, 4213.8, 4217.2, 4220.6, 4224, 4227.4, 
    4230.8, 4234.2, 4237.6, 4241, 4244.4, 4247.8, 4251.2, 4254.6, 4258, 
    4261.4, 4264.8, 4268.2, 4271.6, 4275, 4278.3, 4281.7, 4285.1, 4288.5, 
    4291.9, 4295.2, 4298.6, 4302, 4305.4, 4308.8, 4312.1, 4315.5, 4318.9, 
    4322.3, 4325.7, 4329.1, 4332.5, 4335.8, 4339.2, 4342.6, 4346, 4349.4, 
    4352.9, 4356.3, 4359.7, 4363.1, 4366.5, 4370, 4373.4, 4376.8, 4380.2, 
    4383.6, 4387.1, 4390.5, 4393.9, 4397.3, 4400.8, 4404.2, 4407.6, 4411, 
    4414.4, 4417.9, 4421.3, 4424.7, 4428.1, 4431.6, 4435, 4438.4, 4441.8, 
    4445.3, 4448.7, 4452.1, 4455.6, 4459, 4462.4, 4465.9, 4469.3, 4472.8, 
    4476.2, 4479.6, 4483.1, 4486.5, 4490, 4493.4, 4496.8, 4500.2, 4503.7, 
    4507.1, 4510.5, 4513.9, 4517.3, 4520.7, 4524.1, 4527.6, 4531, 4534.4, 
    4537.8, 4541.2, 4544.6, 4548, 4551.4, 4554.8, 4558.2, 4561.6, 4565.1, 
    4568.5, 4571.9, 4575.3, 4578.7, 4582.1, 4585.4, 4588.8, 4592.2, 4595.6, 
    4599, 4602.3, 4605.7, 4609.1, 4612.4, 4615.8, 4619.1, 4622.5, 4625.9, 
    4629.2, 4632.6, 4636, 4639.4, 4642.7, 4646.1, 4649.5, 4652.9, 4656.3, 
    4659.7, 4663.1, 4666.5, 4669.8, 4673.2, 4676.6, 4680, 4683.5, 4686.9, 
    4690.3, 4693.7, 4697.1, 4700.6, 4704, 4707.4, 4710.8, 4714.3, 4717.7, 
    4721.1, 4724.6, 4728, 4731.4, 4734.9, 4738.3, 4741.7, 4745.2, 4748.6, 
    4752, 4755.5, 4758.9, 4762.3, 4765.8, 4769.2, 4772.7, 4776.1, 4779.5, 
    4783, 4786.4, 4789.9, 4793.3, 4796.7, 4800.2, 4803.6, 4807, 4810.5, 
    4813.9, 4817.3, 4820.8, 4824.2, 4827.6, 4831, 4834.4, 4837.8, 4841.3, 
    4844.7, 4848.1, 4851.5, 4855, 4858.4, 4861.8, 4865.3, 4868.7, 4872.1, 
    4875.6, 4879, 4882.4, 4885.8, 4889.2, 4892.7, 4896.1, 4899.5, 4902.9, 
    4906.3, 4909.7, 4913.1, 4916.5, 4920, 4923.4, 4926.8, 4930.2, 4933.6, 
    4937, 4940.4, 4943.8, 4947.3, 4950.7, 4954.1, 4957.5, 4960.9, 4964.4, 
    4967.8, 4971.2, 4974.6, 4978, 4981.5, 4984.9, 4988.3, 4991.7, 4995.1, 
    4998.5, 5001.9, 5005.4, 5008.8, 5012.2, 5015.6, 5019.1, 5022.5, 5025.9, 
    5029.4, 5032.8, 5036.2, 5039.7, 5043.1, 5046.5, 5049.9, 5053.4, 5056.8, 
    5060.2, 5063.7, 5067.1, 5070.5, 5074, 5077.4, 5080.9, 5084.3, 5087.8, 
    5091.2, 5094.6, 5098, 5101.5, 5104.9, 5108.3, 5111.7, 5115.1, 5118.6, 
    5122, 5125.4, 5128.8, 5132.2, 5135.6, 5139, 5142.4, 5145.8, 5149.2, 
    5152.6, 5156, 5159.4, 5162.8, 5166.2, 5169.6, 5172.9, 5176.3, 5179.7, 
    5183.1, 5186.4, 5189.8, 5193.2, 5196.5, 5199.9, 5203.2, 5206.6, 5209.9, 
    5213.3, 5216.6, 5220, 5223.4, 5226.7, 5230.1, 5233.4, 5236.8, 5240.1, 
    5243.5, 5246.8, 5250.2, 5253.6, 5256.9, 5260.3, 5263.6, 5267, 5270.3, 
    5273.7, 5277.1, 5280.4, 5283.8, 5287.2, 5290.5, 5293.9, 5297.3, 5300.6, 
    5304, 5307.4, 5310.7, 5314.1, 5317.5, 5320.9, 5324.3, 5327.6, 5331, 
    5334.4, 5337.8, 5341.1, 5344.5, 5347.9, 5351.3, 5354.6, 5358, 5361.4, 
    5364.8, 5368.1, 5371.5, 5374.9, 5378.2, 5381.6, 5385, 5388.3, 5391.7, 
    5395.1, 5398.5, 5401.8, 5405.2, 5408.5, 5411.9, 5415.3, 5418.6, 5422, 
    5425.4, 5428.7, 5432.1, 5435.4, 5438.8, 5442.2, 5445.5, 5448.9, 5452.3, 
    5455.6, 5459, 5462.4, 5465.7, 5469.1, 5472.5, 5475.8, 5479.2, 5482.6, 
    5486, 5489.3, 5492.7, 5496.1, 5499.5, 5502.9, 5506.2, 5509.6, 5513, 
    5516.4, 5519.8, 5523.2, 5526.5, 5529.9, 5533.3, 5536.7, 5540.1, 5543.5, 
    5546.8, 5550.2, 5553.6, 5557, 5560.4, 5563.7, 5567.1, 5570.5, 5573.9, 
    5577.2, 5580.6, 5584, 5587.3, 5590.7, 5594, 5597.4, 5600.8, 5604.1, 
    5607.5, 5610.8, 5614.2, 5617.5, 5620.9, 5624.3, 5627.6, 5631, 5634.3, 
    5637.7, 5641.1, 5644.4, 5647.8, 5651.1, 5654.5, 5657.8, 5661.2, 5664.5, 
    5667.9, 5671.2, 5674.5, 5677.9, 5681.2, 5684.6, 5687.9, 5691.3, 5694.6, 
    5698, 5701.3, 5704.7, 5708, 5711.4, 5714.7, 5718.1, 5721.4, 5724.8, 
    5728.1, 5731.5, 5734.9, 5738.2, 5741.6, 5744.9, 5748.2, 5751.6, 5754.9, 
    5758.3, 5761.6, 5765, 5768.3, 5771.6, 5775, 5778.3, 5781.7, 5785, 5788.4, 
    5791.7, 5795.1, 5798.4, 5801.8, 5805.1, 5808.5, 5811.8, 5815.2, 5818.5, 
    5821.9, 5825.2, 5828.6, 5831.9, 5835.3, 5838.6, 5842, 5845.4, 5848.7, 
    5852.1, 5855.4, 5858.7, 5862.1, 5865.4, 5868.8, 5872.1, 5875.5, 5878.8, 
    5882.2, 5885.5, 5888.9, 5892.2, 5895.6, 5898.9, 5902.2, 5905.6, 5908.9, 
    5912.3, 5915.7, 5919, 5922.4, 5925.7, 5929.1, 5932.4, 5935.8, 5939.2, 
    5942.5, 5945.9, 5949.3, 5952.7, 5956, 5959.4, 5962.8, 5966.1, 5969.5, 
    5972.9, 5976.3, 5979.7, 5983, 5986.4, 5989.8, 5993.2, 5996.6, 5999.9, 
    6003.3, 6006.7, 6010.1, 6013.5, 6016.8, 6020.2, 6023.6, 6027, 6030.4, 
    6033.7, 6037.1, 6040.5, 6043.9, 6047.3, 6050.7, 6054.1, 6057.4, 6060.8, 
    6064.2, 6067.6, 6071, 6074.3, 6077.7, 6081.1, 6084.5, 6087.8, 6091.2, 
    6094.6, 6097.9, 6101.3, 6104.6, 6108, 6111.3, 6114.7, 6118, 6121.4, 
    6124.8, 6128.1, 6131.5, 6134.9, 6138.2, 6141.6, 6144.9, 6148.3, 6151.6, 
    6155, 6158.3, 6161.7, 6165, 6168.4, 6171.7, 6175, 6178.4, 6181.7, 6185, 
    6188.4, 6191.7, 6195, 6198.3, 6201.7, 6205, 6208.3, 6211.7, 6215, 6218.3, 
    6221.7, 6225, 6228.4, 6231.7, 6235.1, 6238.4, 6241.7, 6245.1, 6248.4, 
    6251.8, 6255.1, 6258.4, 6261.8, 6265.1, 6268.4, 6271.8, 6275.1, 6278.4, 
    6281.8, 6285.1, 6288.5, 6291.8, 6295.1, 6298.5, 6301.8, 6305.2, 6308.5, 
    6311.9, 6315.2, 6318.6, 6321.9, 6325.3, 6328.6, 6332, 6335.4, 6338.7, 
    6342.1, 6345.4, 6348.8, 6352.1, 6355.4, 6358.8, 6362.1, 6365.5, 6368.8, 
    6372.2, 6375.5, 6378.9, 6382.2, 6385.6, 6389, 6392.4, 6395.7, 6399.1, 
    6402.5, 6405.8, 6409.2, 6412.5, 6415.9, 6419.3, 6422.7, 6426, 6429.4, 
    6432.8, 6436.1, 6439.5, 6442.9, 6446.3, 6449.6, 6453, 6456.4, 6459.8, 
    6463.1, 6466.5, 6469.9, 6473.3, 6476.6, 6480, 6483.4, 6486.8, 6490.1, 
    6493.5, 6496.9, 6500.3, 6503.6, 6507, 6510.4, 6513.8, 6517.1, 6520.5, 
    6523.9, 6527.2, 6530.6, 6534, 6537.4, 6540.7, 6544.1, 6547.5, 6550.8, 
    6554.2, 6557.5, 6560.8, 6564.2, 6567.5, 6570.9, 6574.2, 6577.5, 6580.9, 
    6584.2, 6587.5, 6590.8, 6594.2, 6597.5, 6600.8, 6604.1, 6607.4, 6610.8, 
    6614.1, 6617.4, 6620.7, 6624, 6627.3, 6630.6, 6633.9, 6637.2, 6640.5, 
    6643.8, 6647.1, 6650.4, 6653.7, 6656.9, 6660.2, 6663.5, 6666.8, 6670, 
    6673.3, 6676.6, 6679.9, 6683.1, 6686.4, 6689.7, 6693, 6696.3, 6699.5, 
    6702.8, 6706.1, 6709.4, 6712.7, 6716, 6719.2, 6722.5, 6725.8, 6729.1, 
    6732.4, 6735.7, 6738.9, 6742.2, 6745.5, 6748.8, 6752.1, 6755.4, 6758.7, 
    6762, 6765.3, 6768.6, 6771.9, 6775.2, 6778.5, 6781.8, 6785.1, 6788.4, 
    6791.7, 6795.1, 6798.4, 6801.7, 6805, 6808.3, 6811.6, 6814.9, 6818.2, 
    6821.6, 6824.9, 6828.2, 6831.5, 6834.8, 6838.1, 6841.5, 6844.8, 6848.1, 
    6851.4, 6854.7, 6858.1, 6861.4, 6864.7, 6868, 6871.4, 6874.7, 6878, 
    6881.4, 6884.7, 6888, 6891.4, 6894.7, 6898, 6901.4, 6904.7, 6908, 6911.4, 
    6914.7, 6918, 6921.4, 6924.7, 6928, 6931.4, 6934.7, 6938.1, 6941.4, 
    6944.7, 6948.1, 6951.4, 6954.8, 6958.1, 6961.5, 6964.8, 6968.2, 6971.5, 
    6974.9, 6978.2, 6981.6, 6984.9, 6988.2, 6991.6, 6994.9, 6998.3, 7001.6, 
    7005, 7008.3, 7011.6, 7015, 7018.3, 7021.7, 7025, 7028.4, 7031.7, 7035, 
    7038.4, 7041.7, 7045.1, 7048.4, 7051.8, 7055.1, 7058.5, 7061.8, 7065.2, 
    7068.5, 7071.9, 7075.2, 7078.5, 7081.9, 7085.2, 7088.5, 7091.9, 7095.2, 
    7098.5, 7101.8, 7105.2, 7108.5, 7111.8, 7115.2, 7118.5, 7121.8, 7125.2, 
    7128.5, 7131.8, 7135.2, 7138.5, 7141.8, 7145.2, 7148.5, 7151.8, 7155.2, 
    7158.5, 7161.8, 7165.2, 7168.5, 7171.8, 7175.1, 7178.4, 7181.8, 7185.1, 
    7188.4, 7191.7, 7195, 7198.4, 7201.7, 7205, 7208.3, 7211.7, 7215, 7218.3, 
    7221.6, 7225, 7228.3, 7231.7, 7235, 7238.3, 7241.7, 7245, 7248.3, 7251.7, 
    7255, 7258.4, 7261.7, 7265, 7268.4, 7271.7, 7275, 7278.3, 7281.7, 7285, 
    7288.3, 7291.6, 7295, 7298.3, 7301.6, 7304.9, 7308.3, 7311.6, 7314.9, 
    7318.3, 7321.6, 7324.9, 7328.3, 7331.6, 7334.9, 7338.3, 7341.6, 7344.9, 
    7348.2, 7351.5, 7354.9, 7358.2, 7361.5, 7364.8, 7368.1, 7371.4, 7374.8, 
    7378.1, 7381.4, 7384.7, 7388, 7391.3, 7394.6, 7397.9, 7401.2, 7404.5, 
    7407.9, 7411.2, 7414.5, 7417.8, 7421.1, 7424.4, 7427.7, 7431.1, 7434.4, 
    7437.7, 7441, 7444.3, 7447.6, 7450.9, 7454.2, 7457.5, 7460.8, 7464.1, 
    7467.4, 7470.7, 7474, 7477.3, 7480.6, 7483.9, 7487.3, 7490.6, 7493.9, 
    7497.2, 7500.5, 7503.8, 7507.1, 7510.4, 7513.7, 7517, 7520.3, 7523.6, 
    7526.9, 7530.2, 7533.5, 7536.8, 7540.1, 7543.4, 7546.7, 7550, 7553.3, 
    7556.6, 7559.9, 7563.2, 7566.5, 7569.8, 7573.1, 7576.5, 7579.8, 7583.1, 
    7586.4, 7589.7, 7593, 7596.4, 7599.7, 7603, 7606.3, 7609.6, 7612.9, 
    7616.2, 7619.6, 7622.9, 7626.2, 7629.5, 7632.8, 7636.1, 7639.4, 7642.7, 
    7646, 7649.4, 7652.7, 7656, 7659.3, 7662.6, 7665.9, 7669.2, 7672.6, 
    7675.9, 7679.2, 7682.5, 7685.8, 7689.1, 7692.5, 7695.8, 7699.1, 7702.4, 
    7705.7, 7709, 7712.3, 7715.6, 7718.9, 7722.2, 7725.5, 7728.8, 7732.1, 
    7735.4, 7738.7, 7742, 7745.3, 7748.6, 7751.9, 7755.2, 7758.5, 7761.8, 
    7765.1, 7768.4, 7771.7, 7775, 7778.3, 7781.6, 7784.9, 7788.2, 7791.5, 
    7794.8, 7798.1, 7801.4, 7804.7, 7808, 7811.3, 7814.6, 7817.9, 7821.2, 
    7824.4, 7827.7, 7831, 7834.3, 7837.5, 7840.8, 7844.1, 7847.4, 7850.7, 
    7854, 7857.3, 7860.6, 7863.8, 7867.1, 7870.4, 7873.7, 7877, 7880.3, 
    7883.6, 7886.9, 7890.2, 7893.4, 7896.7, 7900, 7903.3, 7906.5, 7909.8, 
    7913.1, 7916.4, 7919.6, 7922.9, 7926.2, 7929.4, 7932.7, 7936, 7939.2, 
    7942.5, 7945.8, 7949.1, 7952.3, 7955.6, 7958.9, 7962.2, 7965.4, 7968.7, 
    7972, 7975.3, 7978.5, 7981.8, 7985.1, 7988.4, 7991.6, 7994.9, 7998.2, 
    8001.5, 8004.7, 8008, 8011.3, 8014.6, 8017.9, 8021.2, 8024.5, 8027.7, 
    8031, 8034.3, 8037.6, 8040.9, 8044.2, 8047.5, 8050.9, 8054.2, 8057.4, 
    8060.7, 8064, 8067.3, 8070.6, 8073.9, 8077.2, 8080.5, 8083.7, 8087, 
    8090.3, 8093.6, 8096.9, 8100.2, 8103.4, 8106.7, 8110, 8113.3, 8116.6, 
    8119.8, 8123.1, 8126.4, 8129.7, 8132.9, 8136.2, 8139.5, 8142.8, 8146, 
    8149.3, 8152.6, 8155.8, 8159.1, 8162.4, 8165.6, 8168.9, 8172.1, 8175.4, 
    8178.6, 8181.9, 8185.2, 8188.4, 8191.7, 8194.9, 8198.2, 8201.4, 8204.7, 
    8207.9, 8211.2, 8214.5, 8217.8, 8221, 8224.3, 8227.6, 8230.8, 8234.1, 
    8237.4, 8240.7, 8243.9, 8247.2, 8250.5, 8253.8, 8257.1, 8260.3, 8263.6, 
    8266.9, 8270.2, 8273.4, 8276.7, 8280, 8283.3, 8286.6, 8289.9, 8293.1, 
    8296.4, 8299.7, 8303, 8306.3, 8309.6, 8312.9, 8316.2, 8319.5, 8322.8, 
    8326.1, 8329.4, 8332.6, 8335.9, 8339.2, 8342.5, 8345.8, 8349.1, 8352.4, 
    8355.7, 8359, 8362.3, 8365.6, 8368.9, 8372.2, 8375.5, 8378.8, 8382.1, 
    8385.3, 8388.6, 8391.9, 8395.2, 8398.5, 8401.8, 8405, 8408.3, 8411.6, 
    8414.9, 8418.1, 8421.4, 8424.7, 8428, 8431.3, 8434.5, 8437.8, 8441.1, 
    8444.4, 8447.6, 8450.9, 8454.2, 8457.5, 8460.7, 8464, 8467.3, 8470.6, 
    8473.9, 8477.1, 8480.4, 8483.7, 8486.9, 8490.2, 8493.5, 8496.7, 8500, 
    8503.3, 8506.5, 8509.8, 8513.1, 8516.3, 8519.6, 8522.9, 8526.2, 8529.4, 
    8532.7, 8536, 8539.2, 8542.5, 8545.8, 8549, 8552.3, 8555.5, 8558.8, 
    8562.1, 8565.3, 8568.6, 8571.9, 8575.1, 8578.4, 8581.7, 8584.9, 8588.2, 
    8591.4, 8594.7, 8598, 8601.2, 8604.5, 8607.7, 8611, 8614.3, 8617.5, 
    8620.8, 8624.1, 8627.4, 8630.7, 8633.9, 8637.2, 8640.5, 8643.8, 8647.1, 
    8650.4, 8653.6, 8656.9, 8660.2, 8663.5, 8666.8, 8670.1, 8673.3, 8676.6, 
    8679.9, 8683.2, 8686.5, 8689.8, 8693.1, 8696.4, 8699.7, 8702.9, 8706.2, 
    8709.5, 8712.8, 8716.1, 8719.4, 8722.7, 8726, 8729.3, 8732.6, 8735.9, 
    8739.2, 8742.5, 8745.8, 8749.1, 8752.4, 8755.7, 8758.9, 8762.2, 8765.5, 
    8768.8, 8772.1, 8775.3, 8778.6, 8781.9, 8785.2, 8788.5, 8791.8, 8795, 
    8798.3, 8801.6, 8804.9, 8808.2, 8811.5, 8814.8, 8818.1, 8821.4, 8824.6, 
    8827.9, 8831.2, 8834.5, 8837.7, 8841, 8844.3, 8847.5, 8850.8, 8854, 
    8857.3, 8860.5, 8863.8, 8867, 8870.3, 8873.5, 8876.8, 8880, 8883.3, 
    8886.6, 8889.8, 8893.1, 8896.3, 8899.6, 8902.8, 8906.1, 8909.3, 8912.6, 
    8915.8, 8919.1, 8922.3, 8925.5, 8928.8, 8932, 8935.3, 8938.5, 8941.7, 
    8945, 8948.2, 8951.5, 8954.7, 8958, 8961.2, 8964.5, 8967.7, 8971, 8974.2, 
    8977.5, 8980.7, 8984, 8987.2, 8990.4, 8993.7, 8996.9, 9000.2, 9003.4, 
    9006.6, 9009.9, 9013.1, 9016.3, 9019.6, 9022.8, 9026, 9029.3, 9032.5, 
    9035.8, 9039, 9042.2, 9045.5, 9048.7, 9052, 9055.2, 9058.4, 9061.7, 
    9064.9, 9068.2, 9071.4, 9074.6, 9077.9, 9081.1, 9084.3, 9087.6, 9090.8, 
    9094.1, 9097.3, 9100.6, 9103.8, 9107, 9110.3, 9113.5, 9116.8, 9120, 
    9123.3, 9126.5, 9129.8, 9133, 9136.3, 9139.5, 9142.8, 9146, 9149.3, 
    9152.5, 9155.8, 9159, 9162.3, 9165.5, 9168.8, 9172, 9175.3, 9178.5, 
    9181.8, 9185.1, 9188.3, 9191.6, 9194.8, 9198.1, 9201.3, 9204.6, 9207.8, 
    9211.1, 9214.3, 9217.6, 9220.8, 9224.1, 9227.3, 9230.6, 9233.9, 9237.1, 
    9240.4, 9243.7, 9246.9, 9250.2, 9253.5, 9256.7, 9260, 9263.2, 9266.5, 
    9269.8, 9273, 9276.3, 9279.6, 9282.9, 9286.1, 9289.4, 9292.7, 9295.9, 
    9299.2, 9302.5, 9305.8, 9309, 9312.3, 9315.5, 9318.8, 9322.1, 9325.3, 
    9328.6, 9331.9, 9335.1, 9338.4, 9341.6, 9344.9, 9348.1, 9351.4, 9354.7, 
    9357.9, 9361.2, 9364.4, 9367.7, 9370.9, 9374.2, 9377.5, 9380.7, 9384, 
    9387.2, 9390.5, 9393.7, 9397, 9400.2, 9403.5, 9406.7, 9410, 9413.2, 
    9416.5, 9419.7, 9423, 9426.3, 9429.5, 9432.8, 9436, 9439.3, 9442.5, 
    9445.8, 9449.1, 9452.3, 9455.6, 9458.9, 9462.1, 9465.4, 9468.6, 9471.9, 
    9475.2, 9478.4, 9481.7, 9485, 9488.2, 9491.5, 9494.7, 9498, 9501.3, 
    9504.5, 9507.8, 9511, 9514.3, 9517.6, 9520.8, 9524.1, 9527.3, 9530.6, 
    9533.9, 9537.1, 9540.4, 9543.7, 9546.9, 9550.2, 9553.4, 9556.7, 9560, 
    9563.2, 9566.5, 9569.8, 9573, 9576.3, 9579.5, 9582.8, 9586.1, 9589.3, 
    9592.6, 9595.9, 9599.1, 9602.4, 9605.7, 9608.9, 9612.2, 9615.5, 9618.8, 
    9622, 9625.3, 9628.6, 9631.8, 9635.1, 9638.3, 9641.6, 9644.9, 9648.1, 
    9651.4, 9654.6, 9657.9, 9661.1, 9664.3, 9667.6, 9670.8, 9674.1, 9677.3, 
    9680.6, 9683.8, 9687.1, 9690.3, 9693.6, 9696.8, 9700.1, 9703.3, 9706.6, 
    9709.8, 9713.1, 9716.3, 9719.6, 9722.8, 9726.1, 9729.3, 9732.6, 9735.8, 
    9739, 9742.3, 9745.5, 9748.8, 9752, 9755.2, 9758.5, 9761.7, 9764.9, 
    9768.2, 9771.4, 9774.7, 9777.9, 9781.1, 9784.4, 9787.6, 9790.9, 9794.1, 
    9797.4, 9800.6, 9803.8, 9807.1, 9810.3, 9813.5, 9816.8, 9820, 9823.2, 
    9826.5, 9829.7, 9832.9, 9836.2, 9839.4, 9842.6, 9845.9, 9849.1, 9852.4, 
    9855.6, 9858.8, 9862.1, 9865.3, 9868.5, 9871.7, 9875, 9878.2, 9881.4, 
    9884.7, 9887.9, 9891.2, 9894.4, 9897.6, 9900.9, 9904.1, 9907.4, 9910.6, 
    9913.8, 9917.1, 9920.3, 9923.6, 9926.8, 9930.1, 9933.3, 9936.5, 9939.8, 
    9943, 9946.2, 9949.5, 9952.7, 9955.9, 9959.2, 9962.4, 9965.6, 9968.9, 
    9972.1, 9975.4, 9978.6, 9981.8, 9985.1, 9988.3, 9991.6, 9994.8, 9998.1, 
    10001, 10005, 10008, 10011, 10014, 10018, 10021, 10024, 10027, 10031, 
    10034, 10037, 10040, 10043, 10047, 10050, 10053, 10056, 10060, 10063, 
    10066, 10069, 10073, 10076, 10079, 10082, 10086, 10089, 10092, 10095, 
    10098, 10102, 10105, 10108, 10111, 10115, 10118, 10121, 10124, 10128, 
    10131, 10134, 10137, 10140, 10144, 10147, 10150, 10153, 10157, 10160, 
    10163, 10166, 10170, 10173, 10176, 10179, 10183, 10186, 10189, 10192, 
    10195, 10199, 10202, 10205, 10208, 10212, 10215, 10218, 10221, 10225, 
    10228, 10231, 10234, 10238, 10241, 10244, 10247, 10250, 10254, 10257, 
    10260, 10263, 10267, 10270, 10273, 10276, 10279, 10283, 10286, 10289, 
    10292, 10296, 10299, 10302, 10305, 10308, 10312, 10315, 10318, 10321, 
    10324, 10328, 10331, 10334, 10337, 10340, 10344, 10347, 10350, 10353, 
    10357, 10360, 10363, 10366, 10369, 10373, 10376, 10379, 10382, 10386, 
    10389, 10392, 10395, 10399, 10402, 10405, 10408, 10411, 10415, 10418, 
    10421, 10424, 10428, 10431, 10434, 10437, 10441, 10444, 10447, 10450, 
    10454, 10457, 10460, 10463, 10467, 10470, 10473, 10476, 10480, 10483, 
    10486, 10489, 10493, 10496, 10499, 10503, 10506, 10509, 10512, 10516, 
    10519, 10522, 10525, 10529, 10532, 10535, 10538, 10542, 10545, 10548, 
    10552, 10555, 10558, 10561, 10565, 10568, 10571, 10575, 10578, 10581, 
    10584, 10588, 10591, 10594, 10597, 10601, 10604, 10607, 10611, 10614, 
    10617, 10620, 10624, 10627, 10630, 10634, 10637, 10640, 10643, 10647, 
    10650, 10653, 10657, 10660, 10663, 10666, 10670, 10673, 10676, 10680, 
    10683, 10686, 10689, 10693, 10696, 10699, 10703, 10706, 10709, 10712, 
    10716, 10719, 10722, 10726, 10729, 10732, 10736, 10739, 10742, 10745, 
    10749, 10752, 10755, 10759, 10762, 10765, 10769, 10772, 10775, 10778, 
    10782, 10785, 10788, 10792, 10795, 10798, 10802, 10805, 10808, 10812, 
    10815, 10818, 10822, 10825, 10828, 10831, 10835, 10838, 10841, 10845, 
    10848, 10851, 10855, 10858, 10861, 10865, 10868, 10871, 10875, 10878, 
    10881, 10885, 10888, 10891, 10894, 10898, 10901, 10904, 10908, 10911, 
    10914, 10918, 10921, 10924, 10928, 10931, 10934, 10938, 10941, 10944, 
    10948, 10951, 10954, 10958, 10961, 10964, 10968, 10971, 10974, 10978, 
    10981, 10984, 10988, 10991, 10994, 10997, 11001, 11004, 11007, 11011, 
    11014, 11017, 11020, 11024, 11027, 11030, 11033, 11037, 11040, 11043, 
    11046, 11050, 11053, 11056, 11059, 11063, 11066, 11069, 11072, 11075, 
    11079, 11082, 11085, 11088, 11091, 11095, 11098, 11101, 11104, 11107, 
    11111, 11114, 11117, 11120, 11124, 11127, 11130, 11133, 11136, 11140, 
    11143, 11146, 11149, 11153, 11156, 11159, 11162, 11165, 11169, 11172, 
    11175, 11178, 11182, 11185, 11188, 11191, 11194, 11198, 11201, 11204, 
    11207, 11210, 11214, 11217, 11220, 11223, 11227, 11230, 11233, 11236, 
    11239, 11243, 11246, 11249, 11252, 11255, 11259, 11262, 11265, 11268, 
    11271, 11275, 11278, 11281, 11284, 11287, 11291, 11294, 11297, 11300, 
    11304, 11307, 11310, 11313, 11316, 11320, 11323, 11326, 11329, 11333, 
    11336, 11339, 11342, 11346, 11349, 11352, 11355, 11359, 11362, 11365, 
    11368, 11372, 11375, 11378, 11382, 11385, 11388, 11391, 11395, 11398, 
    11401, 11405, 11408, 11411, 11414, 11418, 11421, 11424, 11427, 11431, 
    11434, 11437, 11441, 11444, 11447, 11450, 11454, 11457, 11460, 11463, 
    11467, 11470, 11473, 11477, 11480, 11483, 11486, 11490, 11493, 11496, 
    11499, 11503, 11506, 11509, 11512, 11516, 11519, 11522, 11525, 11529, 
    11532, 11535, 11539, 11542, 11545, 11548, 11552, 11555, 11558, 11562, 
    11565, 11568, 11571, 11575, 11578, 11581, 11585, 11588, 11591, 11594, 
    11598, 11601, 11604, 11607, 11611, 11614, 11617, 11621, 11624, 11627, 
    11630, 11634, 11637, 11640, 11643, 11647, 11650, 11653, 11656, 11660, 
    11663, 11666, 11669, 11672, 11676, 11679, 11682, 11685, 11689, 11692, 
    11695, 11698, 11702, 11705, 11708, 11711, 11715, 11718, 11721, 11725, 
    11728, 11731, 11734, 11738, 11741, 11744, 11748, 11751, 11754, 11757, 
    11761, 11764, 11767, 11770, 11774, 11777, 11780, 11784, 11787, 11790, 
    11793, 11797, 11800, 11803, 11807, 11810, 11813, 11816, 11820, 11823, 
    11826, 11829, 11833, 11836, 11839, 11842, 11846, 11849, 11852, 11855, 
    11859, 11862, 11865, 11869, 11872, 11875, 11878, 11882, 11885, 11888, 
    11891, 11895, 11898, 11901, 11904, 11908, 11911, 11914, 11918, 11921, 
    11924, 11927, 11931, 11934, 11937, 11941, 11944, 11947, 11950, 11954, 
    11957, 11960, 11963, 11967, 11970, 11973, 11976, 11980, 11983, 11986, 
    11989, 11993, 11996, 11999, 12002, 12006, 12009, 12012, 12015, 12019, 
    12022, 12025, 12028, 12032, 12035, 12038, 12041, 12045, 12048, 12051, 
    12054, 12058, 12061, 12064, 12067, 12071, 12074, 12077, 12080, 12084, 
    12087, 12090, 12093, 12096, 12100, 12103, 12106, 12109, 12113, 12116, 
    12119, 12122, 12125, 12129, 12132, 12135, 12138, 12141, 12145, 12148, 
    12151, 12154, 12157, 12161, 12164, 12167, 12170, 12173, 12177, 12180, 
    12183, 12186, 12189, 12193, 12196, 12199, 12202, 12205, 12209, 12212, 
    12215, 12218, 12221, 12225, 12228, 12231, 12234, 12238, 12241, 12244, 
    12247, 12250, 12254, 12257, 12260, 12263, 12267, 12270, 12273, 12276, 
    12280, 12283, 12286, 12289, 12292, 12296, 12299, 12302, 12305, 12309, 
    12312, 12315, 12318, 12322, 12325, 12328, 12331, 12335, 12338, 12341, 
    12344, 12347, 12351, 12354, 12357, 12360, 12364, 12367, 12370, 12373, 
    12376, 12380, 12383, 12386, 12389, 12393, 12396, 12399, 12402, 12406, 
    12409, 12412, 12415, 12419, 12422, 12425, 12428, 12431, 12435, 12438, 
    12441, 12444, 12448, 12451, 12454, 12457, 12461, 12464, 12467, 12470, 
    12473, 12477, 12480, 12483, 12486, 12489, 12493, 12496, 12499, 12502, 
    12505, 12509, 12512, 12515, 12518, 12521, 12525, 12528, 12531, 12534, 
    12537, 12541, 12544, 12547, 12550, 12553, 12557, 12560, 12563, 12566, 
    12569, 12573, 12576, 12579, 12582, 12585, 12589, 12592, 12595, 12598, 
    12601, 12605, 12608, 12611, 12614, 12617, 12621, 12624, 12627, 12630, 
    12633, 12637, 12640, 12643, 12646, 12650, 12653, 12656, 12659, 12662, 
    12666, 12669, 12672, 12675, 12678, 12682, 12685, 12688, 12691, 12694, 
    12698, 12701, 12704, 12707, 12711, 12714, 12717, 12720, 12723, 12727, 
    12730, 12733, 12736, 12739, 12743, 12746, 12749, 12752, 12755, 12759, 
    12762, 12765, 12768, 12771, 12775, 12778, 12781, 12784, 12787, 12791, 
    12794, 12797, 12800, 12803, 12806, 12810, 12813, 12816, 12819, 12822, 
    12825, 12829, 12832, 12835, 12838, 12841, 12845, 12848, 12851, 12854, 
    12857, 12860, 12864, 12867, 12870, 12873, 12876, 12879, 12883, 12886, 
    12896, 12907, 12917, 12927, 12937, 12947, 12957, 12966, 12976, 12985, 
    12995, 13004, 13014, 13024, 13034, 13044, 13055, 13066, 13077, 13088, 
    13100, 13112, 13124, 13136, 13149, 13162, 13175, 13188, 13201, 13214, 
    13228, 13241, 13254, 13267, 13280, 13292, 13305, 13317, 13329, 13341, 
    13353, 13365, 13377, 13388, 13400, 13411, 13423, 13434, 13446, 13457, 
    13469, 13480, 13492, 13504, 13516, 13528, 13540, 13552, 13565, 13577, 
    13590, 13602, 13615, 13628, 13640, 13653, 13666, 13679, 13691, 13704, 
    13717, 13729, 13742, 13754, 13767, 13779, 13791, 13803, 13816, 13828, 
    13840, 13852, 13864, 13877, 13889, 13901, 13914, 13926, 13939, 13951, 
    13964, 13977, 13990, 14003, 14016, 14029, 14043, 14056, 14069, 14083, 
    14096, 14110, 14123, 14137, 14150, 14164, 14178, 14191, 14205, 14218, 
    14232, 14246, 14259, 14273, 14286, 14300, 14313, 14327, 14340, 14354, 
    14367, 14380, 14394, 14407, 14420, 14433, 14446, 14460, 14473, 14486, 
    14499, 14512, 14525, 14538, 14551, 14564, 14577, 14590, 14603, 14616, 
    14629, 14642, 14656, 14669, 14683, 14696, 14710, 14724, 14738, 14752, 
    14766, 14780, 14795, 14810, 14824, 14839, 14854, 14870, 14885, 14900, 
    14916, 14931, 14947, 14962, 14978, 14994, 15010, 15025, 15041, 15057, 
    15073, 15089, 15104, 15120, 15136, 15152, 15167, 15183, 15199, 15214, 
    15230, 15246, 15261, 15277, 15293, 15308, 15324, 15339, 15355, 15371, 
    15386, 15402, 15418, 15433, 15449, 15464, 15480, 15496, 15512, 15527, 
    15543, 15559, 15575, 15591, 15607, 15624, 15640, 15657, 15674, 15691, 
    15709, 15727, 15745, 15763, 15781, 15800, 15819, 15838, 15858, 15878, 
    15898, 15918, 15938, 15958, 15979, 16000, 16020, 16041, 16062, 16082, 
    16103, 16124, 16145, 16165, 16186, 16207, 16227, 16248, 16268, 16289, 
    16309, 16329, 16350, 16370, 16390, 16410, 16431, 16451, 16471, 16490, 
    16510, 16530, 16549, 16568, 16588, 16607, 16625, 16644, 16662, 16680, 
    16698, 16715, 16732, 16749, 16766, 16783, 16799, 16815, 16831, 16847, 
    16862, 16877, 16893, 16908, 16923, 16938, 16953, 16968, 16983, 16998, 
    17013, 17028, 17043, 17059, 17074, 17089, 17105, 17120, 17136, 17151, 
    17167, 17183, 17198, 17214, 17229, 17245, 17261, 17277, 17292, 17308, 
    17324, 17341, 17357, 17373, 17390, 17407, 17424, 17441, 17459, 17476, 
    17494, 17512, 17531, 17550, 17569, 17588, 17607, 17627, 17647, 17667, 
    17687, 17707, 17728, 17749, 17770, 17791, 17813, 17835, 17856, 17878, 
    17900, 17922, 17945, 17967, 17990, 18012, 18035, 18057, 18080, 18103, 
    18126, 18148, 18171, 18194, 18216, 18239, 18261, 18284, 18306, 18328, 
    18351, 18373, 18395, 18416, 18438, 18460, 18481, 18503, 18524, 18545, 
    18566, 18587, 18608, 18629, 18650, 18670, 18690, 18711, 18731, 18751, 
    18771, 18791, 18811, 18831, 18850, 18870, 18890, 18909, 18929, 18948, 
    18968, 18987, 19007, 19026, 19045, 19065, 19084, 19103, 19123, 19142, 
    19161, 19180, 19200, 19219, 19238, 19257, 19277, 19296, 19315, 19335, 
    19354, 19374, 19394, 19413, 19433, 19454, 19474, 19494, 19515, 19536, 
    19557, 19578, 19600, 19621, 19643, 19665, 19687, 19709, 19731, 19753, 
    19775, 19797, 19820, 19842, 19864, 19886, 19908, 19930, 19952, 19974, 
    19995, 20017, 20039, 20060, 20082, 20103, 20125, 20146, 20168, 20190, 
    20211, 20233, 20255, 20276, 20298, 20320, 20342, 20364, 20386, 20409, 
    20431, 20453, 20475, 20498, 20520, 20543, 20565, 20588, 20610, 20633, 
    20656, 20679, 20702, 20726, 20749, 20773, 20797, 20821, 20846, 20870, 
    20895, 20920, 20945, 20970, 20996, 21022, 21047, 21073, 21099, 21125, 
    21152, 21178, 21204, 21230, 21256, 21282, 21308, 21334, 21360, 21385, 
    21411, 21436, 21461, 21486, 21511, 21535, 21560, 21584, 21607, 21631, 
    21654, 21678, 21701, 21723, 21746, 21769, 21791, 21813, 21836, 21858, 
    21880, 21902, 21925, 21947, 21970, 21992, 22015, 22038, 22062, 22085, 
    22109, 22133, 22158, 22182, 22207, 22233, 22259, 22284, 22311, 22337, 
    22364, 22391, 22418, 22445, 22473, 22500, 22528, 22556, 22584, 22611, 
    22639, 22667, 22695, 22723, 22751, 22778, 22806, 22834, 22861, 22889, 
    22916, 22944, 22971, 22999, 23026, 23053, 23081, 23108, 23136, 23163, 
    23190, 23217, 23245, 23272, 23299, 23326, 23353, 23379, 23406, 23432, 
    23459, 23485, 23511, 23536, 23562, 23587, 23613, 23638, 23663, 23688, 
    23713, 23738, 23763, 23787, 23812, 23837, 23862, 23887, 23912, 23938, 
    23963, 23989, 24015, 24041, 24067, 24093, 24120, 24147, 24174, 24201, 
    24228, 24256, 24284, 24312, 24341, 24369, 24398, 24427, 24456, 24486, 
    24515, 24545, 24575, 24605, 24635, 24666, 24696, 24726, 24757, 24787, 
    24818, 24848, 24879, 24909, 24940, 24970, 25000, 25031, 25061, 25091, 
    25121, 25151, 25182, 25212, 25242, 25271, 25301, 25331, 25361, 25391, 
    25420, 25450, 25480, 25509, 25539, 25568, 25597, 25627, 25656, 25685, 
    25715, 25744, 25773, 25802, 25832, 25861, 25890, 25919, 25949, 25978, 
    26007, 26036, 26065, 26094, 26123, 26152, 26181, 26209, 26238, 26266, 
    26294, 26323, 26351, 26379, 26407, 26435, 26463, 26491, 26519, 26547, 
    26576, 26605, 26633, 26662, 26691, 26721, 26750, 26780, 26810, 26840, 
    26871, 26902, 26933, 26964, 26995, 27027, 27059, 27091, 27124, 27156, 
    27189, 27222, 27255, 27288, 27322, 27355, 27389, 27423, 27456, 27490, 
    27523, 27557, 27590, 27624, 27657, 27691, 27724, 27757, 27790, 27823, 
    27855, 27888, 27921, 27953, 27985, 28018, 28050, 28082, 28114, 28146, 
    28178, 28210, 28242, 28274, 28306, 28337, 28369, 28401, 28433, 28465, 
    28496, 28528, 28560, 28592, 28624, 28655, 28687, 28719, 28751, 28783, 
    28815, 28846, 28878, 28910, 28942, 28974, 29006, 29037, 29069, 29101, 
    29133, 29165, 29196, 29228, 29260, 29291, 29323, 29354, 29386, 29417, 
    29448, 29480, 29511, 29542, 29574, 29605, 29636, 29667, 29698, 29729, 
    29760, 29792, 29823, 29854, 29886, 29918, 29949, 29981, 30013, 30046, 
    30078, 30111, 30143, 30176, 30209, 30243, 30276, 30310, 30343, 30377, 
    30411, 30445, 30479, 30514, 30548, 30582, 30617, 30651, 30685, 30720, 
    30754, 30788, 30822, 30857, 30891, 30925, 30959, 30993, 31027, 31061, 
    31095, 31129, 31163, 31197, 31231, 31265, 31298, 31332, 31366, 31400, 
    31434, 31468, 31502, 31536, 31570, 31604, 31638, 31672, 31706, 31741, 
    31775, 31810, 31844, 31879, 31914, 31948, 31983, 32018, 32053, 32088, 
    32123, 32158, 32193, 32228, 32262, 32297, 32332, 32367, 32402, 32437, 
    32471, 32506, 32541, 32576, 32611, 32645, 32680, 32715, 32750, 32785, 
    32820, 32855, 32890, 32925, 32960, 32996, 33031, 33066, 33101, 33137, 
    33172, 33207, 33243, 33278, 33313, 33349, 33384, 33419, 33455, 33490, 
    33525, 33560, 33595, 33630, 33665, 33700, 33735, 33770, 33805, 33840, 
    33874, 33909, 33944, 33978, 34013, 34048, 34082, 34117, 34151, 34186, 
    34221, 34255, 34290, 34324, 34359, 34394, 34428, 34463, 34498, 34532, 
    34567, 34602, 34637, 34671, 34706, 34741, 34776, 34811, 34846, 34882, 
    34917, 34952, 34988, 35023, 35059, 35094, 35130, 35166, 35201, 35237, 
    35273, 35309, 35344, 35380, 35416, 35451, 35487, 35522, 35557, 35593, 
    35628, 35663, 35698, 35734, 35769, 35804, 35839, 35874, 35910, 35945, 
    35980, 36016, 36051, 36087, 36123, 36158, 36194, 36230, 36266, 36302, 
    36338, 36374, 36411, 36447, 36483, 36519, 36555, 36592, 36628, 36664, 
    36700, 36736, 36772, 36808, 36844, 36880, 36916, 36951, 36987, 37022, 
    37058, 37093, 37129, 37164, 37199, 37234, 37269, 37304, 37339, 37374, 
    37409, 37444, 37479, 37513, 37548, 37583, 37618, 37653, 37688, 37723, 
    37758, 37794, 37829, 37864, 37900, 37935, 37971, 38007, 38043, 38079, 
    38115, 38151, 38187, 38224, 38260, 38297, 38334, 38370, 38407, 38444, 
    38481, 38518, 38555, 38592, 38629, 38666, 38703, 38740, 38776, 38813, 
    38850, 38887, 38924, 38960, 38997, 39034, 39070, 39107, 39143, 39180, 
    39216, 39252, 39288, 39325, 39361, 39397, 39433, 39469, 39506, 39542, 
    39578, 39614, 39650, 39686, 39722, 39757, 39793, 39829, 39865, 39901, 
    39937, 39973, 40008, 40044, 40080, 40116, 40152, 40188, 40224, 40260, 
    40296, 40331, 40367, 40403, 40439, 40475, 40511, 40548, 40584, 40620, 
    40656, 40692, 40728, 40764, 40800, 40836, 40872, 40909, 40945, 40981, 
    41017, 41053, 41090, 41126, 41162, 41199, 41235, 41271, 41308, 41344, 
    41381, 41417, 41454, 41490, 41527, 41563, 41599, 41636, 41672, 41709, 
    41745, 41782, 41818, 41855, 41891, 41928, 41964, 42000, 42037, 42073, 
    42110, 42146, 42182, 42219, 42255, 42291, 42328, 42364, 42400, 42437, 
    42473, 42509, 42546, 42582, 42618, 42655, 42691, 42727, 42764, 42800, 
    42837, 42873, 42910, 42946, 42983, 43020, 43056, 43093, 43130, 43167, 
    43204, 43241, 43277, 43314, 43351, 43388, 43425, 43462, 43499, 43536, 
    43573, 43610, 43647, 43684, 43721, 43758, 43794, 43831, 43868, 43905, 
    43942, 43979, 44015, 44052, 44089, 44125, 44162, 44199, 44235, 44272, 
    44308, 44345, 44381, 44418, 44455, 44492, 44528, 44565, 44602, 44639, 
    44676, 44713, 44751, 44788, 44825, 44863, 44900, 44938, 44975, 45012, 
    45050, 45087, 45125, 45162, 45199, 45236, 45273, 45309, 45346, 45382, 
    45418, 45454, 45490, 45526, 45561, 45597, 45632, 45667, 45702, 45737, 
    45772, 45807, 45842, 45877, 45913, 45948, 45983, 46019, 46054, 46090, 
    46126, 46162, 46198, 46234, 46270, 46307, 46344, 46381, 46418, 46455, 
    46492, 46529, 46567, 46604, 46642, 46680, 46717, 46755, 46793, 46830, 
    46868, 46905, 46943, 46980, 47018, 47055, 47092, 47130, 47167, 47203, 
    47240, 47277, 47313, 47350, 47386, 47422, 47458, 47494, 47530, 47566, 
    47601, 47637, 47673, 47708, 47744, 47779, 47815, 47851, 47886, 47922, 
    47958, 47993, 48029, 48065, 48100, 48136, 48172, 48208, 48244, 48280, 
    48316, 48352, 48388, 48424, 48460, 48496, 48532, 48569, 48605, 48641, 
    48678, 48714, 48751, 48787, 48824, 48861, 48898, 48935, 48972, 49009, 
    49046, 49084, 49121, 49159, 49196, 49234, 49271, 49309, 49346, 49383, 
    49421, 49458, 49496, 49533, 49570, 49607, 49644, 49681, 49718, 49755, 
    49792, 49829, 49866, 49903, 49939, 49976, 50013, 50050, 50086, 50123, 
    50160, 50196, 50233, 50270, 50306, 50343, 50379, 50416, 50453, 50489, 
    50525, 50562, 50598, 50634, 50671, 50707, 50743, 50779, 50815, 50851, 
    50887, 50923, 50959, 50994, 51030, 51066, 51102, 51138, 51174, 51210, 
    51246, 51282, 51318, 51354, 51390, 51426, 51462, 51498, 51534, 51570, 
    51606, 51642, 51678, 51714, 51749, 51785, 51821, 51856, 51892, 51927, 
    51963, 51998, 52034, 52069, 52105, 52140, 52176, 52212, 52247, 52283, 
    52319, 52354, 52390, 52426, 52462, 52498, 52534, 52569, 52605, 52641, 
    52677, 52713, 52749, 52786, 52822, 52858, 52894, 52930, 52966, 53003, 
    53039, 53076, 53112, 53149, 53185, 53222, 53259, 53295, 53332, 53369, 
    53405, 53442, 53479, 53515, 53552, 53588, 53625, 53661, 53698, 53734, 
    53770, 53806, 53843, 53879, 53915, 53951, 53987, 54023, 54060, 54096, 
    54132, 54168, 54204, 54240, 54277, 54313, 54349, 54385, 54422, 54458, 
    54494, 54531, 54567, 54603, 54640, 54676, 54712, 54749, 54785, 54821, 
    54858, 54894, 54930, 54967, 55003, 55039, 55076, 55112, 55148, 55185, 
    55221, 55257, 55293, 55330, 55366, 55402, 55438, 55475, 55511, 55547, 
    55583, 55619, 55655, 55691, 55727, 55763, 55799, 55835, 55871, 55907, 
    55943, 55979, 56015, 56051, 56087, 56123, 56159, 56195, 56231, 56268, 
    56304, 56341, 56377, 56414, 56451, 56488, 56524, 56561, 56599, 56636, 
    56673, 56710, 56747, 56784, 56821, 56858, 56895, 56932, 56969, 57006, 
    57043, 57079, 57116, 57152, 57188, 57225, 57261, 57297, 57333, 57369, 
    57405, 57441, 57476, 57512, 57548, 57584, 57620, 57656, 57691, 57727, 
    57763, 57799, 57835, 57871, 57907, 57943, 57979, 58015, 58051, 58087, 
    58122, 58158, 58194, 58230, 58266, 58302, 58338, 58374, 58410, 58446, 
    58482, 58518, 58554, 58590, 58626, 58662, 58699, 58735, 58771, 58807, 
    58843, 58879, 58916, 58952, 58988, 59025, 59061, 59097, 59134, 59170, 
    59207, 59244, 59280, 59317, 59353, 59390, 59427, 59463 ;

 refrac =
  296.3, 296.54, 296.78, 297.03, 297.29, 297.55, 297.8, 298.05, 298.29, 
    298.53, 298.76, 298.98, 299.18, 299.37, 299.54, 299.69, 299.82, 299.93, 
    300.02, 300.08, 300.13, 300.16, 300.17, 300.17, 300.16, 300.15, 300.13, 
    300.1, 300.06, 300.02, 299.97, 299.93, 299.87, 299.81, 299.74, 299.66, 
    299.56, 299.46, 299.35, 299.23, 299.1, 298.97, 298.84, 298.69, 298.54, 
    298.39, 298.25, 298.1, 297.96, 297.81, 297.67, 297.53, 297.39, 297.26, 
    297.12, 296.99, 296.86, 296.74, 296.62, 296.5, 296.38, 296.25, 296.12, 
    295.98, 295.84, 295.7, 295.56, 295.43, 295.3, 295.16, 295.03, 294.89, 
    294.77, 294.64, 294.52, 294.41, 294.3, 294.19, 294.08, 293.98, 293.87, 
    293.77, 293.68, 293.58, 293.48, 293.38, 293.27, 293.16, 293.05, 292.94, 
    292.82, 292.71, 292.59, 292.47, 292.35, 292.22, 292.09, 291.96, 291.82, 
    291.69, 291.55, 291.42, 291.28, 291.14, 291, 290.86, 290.72, 290.58, 
    290.44, 290.29, 290.15, 290, 289.86, 289.71, 289.56, 289.41, 289.27, 
    289.12, 288.97, 288.83, 288.68, 288.54, 288.41, 288.27, 288.14, 288, 
    287.87, 287.75, 287.62, 287.49, 287.37, 287.24, 287.12, 286.99, 286.87, 
    286.74, 286.61, 286.49, 286.36, 286.23, 286.1, 285.97, 285.84, 285.71, 
    285.58, 285.45, 285.32, 285.19, 285.06, 284.93, 284.79, 284.66, 284.53, 
    284.41, 284.28, 284.14, 284.01, 283.87, 283.74, 283.6, 283.45, 283.3, 
    283.15, 282.99, 282.83, 282.67, 282.5, 282.33, 282.15, 281.98, 281.79, 
    281.61, 281.42, 281.22, 281.03, 280.83, 280.63, 280.42, 280.21, 280, 
    279.77, 279.55, 279.31, 279.07, 278.82, 278.55, 278.28, 277.98, 277.68, 
    277.36, 277.02, 276.66, 276.3, 275.92, 275.55, 275.18, 274.81, 274.44, 
    274.07, 273.71, 273.35, 273, 272.65, 272.3, 271.95, 271.6, 271.25, 270.9, 
    270.54, 270.18, 269.83, 269.48, 269.13, 268.77, 268.42, 268.08, 267.75, 
    267.43, 267.11, 266.81, 266.5, 266.21, 265.92, 265.65, 265.38, 265.14, 
    264.91, 264.69, 264.5, 264.32, 264.15, 263.99, 263.83, 263.68, 263.52, 
    263.35, 263.19, 263.02, 262.84, 262.65, 262.46, 262.28, 262.1, 261.92, 
    261.75, 261.58, 261.42, 261.26, 261.11, 260.96, 260.81, 260.68, 260.56, 
    260.44, 260.31, 260.18, 260.05, 259.91, 259.79, 259.66, 259.54, 259.43, 
    259.33, 259.23, 259.13, 259.03, 258.94, 258.85, 258.77, 258.7, 258.62, 
    258.55, 258.49, 258.43, 258.37, 258.32, 258.28, 258.24, 258.21, 258.19, 
    258.16, 258.14, 258.11, 258.09, 258.08, 258.06, 258.05, 258.03, 258.01, 
    257.99, 257.96, 257.92, 257.89, 257.86, 257.83, 257.8, 257.77, 257.74, 
    257.71, 257.67, 257.62, 257.56, 257.5, 257.44, 257.37, 257.3, 257.22, 
    257.15, 257.07, 256.99, 256.91, 256.83, 256.75, 256.68, 256.6, 256.52, 
    256.45, 256.38, 256.3, 256.23, 256.16, 256.09, 256.02, 255.94, 255.86, 
    255.77, 255.69, 255.6, 255.51, 255.43, 255.35, 255.27, 255.2, 255.13, 
    255.06, 255, 254.94, 254.89, 254.84, 254.8, 254.77, 254.74, 254.72, 
    254.7, 254.68, 254.66, 254.64, 254.62, 254.6, 254.57, 254.54, 254.51, 
    254.47, 254.44, 254.39, 254.35, 254.3, 254.25, 254.2, 254.15, 254.11, 
    254.06, 254.02, 253.98, 253.94, 253.9, 253.86, 253.83, 253.78, 253.73, 
    253.68, 253.63, 253.57, 253.51, 253.44, 253.37, 253.3, 253.22, 253.14, 
    253.05, 252.96, 252.87, 252.78, 252.68, 252.59, 252.5, 252.4, 252.31, 
    252.21, 252.12, 252.03, 251.93, 251.84, 251.74, 251.64, 251.54, 251.44, 
    251.33, 251.23, 251.13, 251.02, 250.92, 250.82, 250.72, 250.63, 250.53, 
    250.43, 250.34, 250.25, 250.15, 250.06, 249.97, 249.89, 249.8, 249.71, 
    249.63, 249.54, 249.45, 249.36, 249.27, 249.18, 249.1, 249.01, 248.92, 
    248.83, 248.75, 248.66, 248.58, 248.49, 248.41, 248.33, 248.25, 248.17, 
    248.09, 248.01, 247.93, 247.85, 247.77, 247.69, 247.61, 247.52, 247.43, 
    247.34, 247.25, 247.17, 247.08, 246.99, 246.9, 246.81, 246.72, 246.64, 
    246.55, 246.46, 246.37, 246.29, 246.21, 246.12, 246.04, 245.96, 245.87, 
    245.79, 245.71, 245.63, 245.55, 245.46, 245.37, 245.29, 245.2, 245.11, 
    245.03, 244.95, 244.86, 244.78, 244.7, 244.62, 244.54, 244.47, 244.39, 
    244.32, 244.25, 244.18, 244.11, 244.04, 243.97, 243.9, 243.82, 243.74, 
    243.67, 243.58, 243.5, 243.41, 243.33, 243.24, 243.15, 243.06, 242.97, 
    242.88, 242.79, 242.7, 242.61, 242.52, 242.43, 242.34, 242.25, 242.16, 
    242.07, 241.99, 241.9, 241.81, 241.71, 241.62, 241.53, 241.44, 241.34, 
    241.25, 241.15, 241.05, 240.95, 240.85, 240.75, 240.65, 240.55, 240.46, 
    240.36, 240.26, 240.16, 240.06, 239.97, 239.87, 239.77, 239.68, 239.58, 
    239.48, 239.39, 239.29, 239.19, 239.1, 239, 238.9, 238.8, 238.7, 238.6, 
    238.5, 238.41, 238.31, 238.21, 238.11, 238.02, 237.92, 237.82, 237.73, 
    237.63, 237.53, 237.44, 237.34, 237.25, 237.15, 237.06, 236.97, 236.87, 
    236.78, 236.69, 236.59, 236.5, 236.41, 236.32, 236.23, 236.14, 236.05, 
    235.96, 235.86, 235.77, 235.68, 235.58, 235.49, 235.39, 235.3, 235.2, 
    235.1, 235, 234.9, 234.79, 234.69, 234.59, 234.48, 234.38, 234.27, 
    234.16, 234.06, 233.95, 233.85, 233.74, 233.63, 233.53, 233.42, 233.32, 
    233.21, 233.1, 233, 232.89, 232.78, 232.68, 232.57, 232.46, 232.35, 
    232.24, 232.13, 232.03, 231.92, 231.81, 231.71, 231.61, 231.51, 231.41, 
    231.31, 231.21, 231.12, 231.03, 230.94, 230.85, 230.76, 230.66, 230.57, 
    230.49, 230.4, 230.31, 230.22, 230.13, 230.05, 229.96, 229.87, 229.78, 
    229.69, 229.6, 229.5, 229.41, 229.32, 229.22, 229.13, 229.04, 228.94, 
    228.85, 228.76, 228.67, 228.59, 228.5, 228.41, 228.33, 228.24, 228.16, 
    228.07, 227.99, 227.91, 227.82, 227.74, 227.66, 227.57, 227.49, 227.41, 
    227.33, 227.25, 227.16, 227.08, 227, 226.92, 226.83, 226.75, 226.67, 
    226.59, 226.5, 226.42, 226.34, 226.26, 226.18, 226.1, 226.03, 225.95, 
    225.88, 225.81, 225.73, 225.66, 225.59, 225.51, 225.44, 225.36, 225.28, 
    225.2, 225.12, 225.04, 224.95, 224.86, 224.77, 224.68, 224.59, 224.49, 
    224.39, 224.29, 224.19, 224.09, 223.99, 223.89, 223.78, 223.67, 223.57, 
    223.46, 223.36, 223.25, 223.15, 223.04, 222.94, 222.84, 222.74, 222.64, 
    222.53, 222.43, 222.33, 222.23, 222.13, 222.02, 221.92, 221.82, 221.72, 
    221.62, 221.52, 221.42, 221.32, 221.22, 221.12, 221.03, 220.93, 220.84, 
    220.74, 220.65, 220.56, 220.47, 220.38, 220.29, 220.2, 220.12, 220.03, 
    219.94, 219.86, 219.78, 219.7, 219.61, 219.53, 219.45, 219.37, 219.28, 
    219.2, 219.12, 219.04, 218.96, 218.88, 218.79, 218.71, 218.63, 218.55, 
    218.47, 218.39, 218.31, 218.23, 218.15, 218.07, 218, 217.92, 217.84, 
    217.76, 217.68, 217.6, 217.51, 217.42, 217.33, 217.23, 217.12, 217.02, 
    216.91, 216.8, 216.69, 216.57, 216.45, 216.33, 216.2, 216.07, 215.94, 
    215.81, 215.67, 215.53, 215.39, 215.25, 215.1, 214.95, 214.79, 214.64, 
    214.48, 214.31, 214.15, 213.98, 213.81, 213.63, 213.45, 213.27, 213.08, 
    212.89, 212.7, 212.5, 212.31, 212.11, 211.9, 211.7, 211.5, 211.3, 211.09, 
    210.89, 210.69, 210.48, 210.28, 210.07, 209.87, 209.67, 209.46, 209.26, 
    209.06, 208.85, 208.65, 208.45, 208.24, 208.04, 207.84, 207.65, 207.45, 
    207.26, 207.07, 206.88, 206.69, 206.51, 206.33, 206.15, 205.98, 205.81, 
    205.64, 205.48, 205.32, 205.16, 205.01, 204.87, 204.72, 204.59, 204.46, 
    204.33, 204.2, 204.09, 203.97, 203.86, 203.75, 203.65, 203.54, 203.44, 
    203.34, 203.24, 203.15, 203.05, 202.96, 202.87, 202.78, 202.7, 202.61, 
    202.53, 202.44, 202.36, 202.28, 202.2, 202.11, 202.03, 201.95, 201.86, 
    201.78, 201.7, 201.61, 201.52, 201.44, 201.35, 201.26, 201.17, 201.09, 
    201, 200.91, 200.82, 200.73, 200.64, 200.55, 200.46, 200.37, 200.28, 
    200.19, 200.11, 200.02, 199.93, 199.84, 199.76, 199.67, 199.59, 199.5, 
    199.42, 199.33, 199.25, 199.16, 199.08, 199, 198.91, 198.83, 198.74, 
    198.66, 198.58, 198.49, 198.41, 198.33, 198.25, 198.17, 198.09, 198.01, 
    197.93, 197.85, 197.78, 197.7, 197.63, 197.55, 197.48, 197.41, 197.34, 
    197.27, 197.2, 197.13, 197.06, 197, 196.93, 196.86, 196.79, 196.72, 
    196.66, 196.59, 196.52, 196.45, 196.39, 196.32, 196.25, 196.19, 196.12, 
    196.05, 195.99, 195.92, 195.86, 195.79, 195.73, 195.67, 195.6, 195.54, 
    195.48, 195.41, 195.35, 195.29, 195.22, 195.16, 195.09, 195.02, 194.95, 
    194.89, 194.82, 194.76, 194.69, 194.62, 194.56, 194.49, 194.43, 194.37, 
    194.31, 194.25, 194.18, 194.12, 194.06, 194, 193.94, 193.87, 193.81, 
    193.75, 193.69, 193.62, 193.56, 193.49, 193.43, 193.36, 193.3, 193.23, 
    193.17, 193.1, 193.04, 192.97, 192.9, 192.84, 192.77, 192.71, 192.64, 
    192.57, 192.51, 192.44, 192.37, 192.3, 192.23, 192.16, 192.09, 192.02, 
    191.95, 191.88, 191.8, 191.73, 191.65, 191.58, 191.5, 191.42, 191.35, 
    191.27, 191.19, 191.11, 191.03, 190.95, 190.87, 190.79, 190.71, 190.64, 
    190.56, 190.48, 190.4, 190.32, 190.25, 190.17, 190.1, 190.02, 189.95, 
    189.87, 189.8, 189.72, 189.65, 189.57, 189.5, 189.43, 189.35, 189.28, 
    189.2, 189.13, 189.05, 188.98, 188.9, 188.83, 188.76, 188.69, 188.61, 
    188.54, 188.47, 188.4, 188.34, 188.27, 188.2, 188.14, 188.07, 188.01, 
    187.94, 187.88, 187.81, 187.75, 187.68, 187.62, 187.55, 187.48, 187.41, 
    187.35, 187.28, 187.21, 187.15, 187.08, 187.01, 186.95, 186.88, 186.81, 
    186.75, 186.68, 186.62, 186.55, 186.49, 186.42, 186.36, 186.29, 186.23, 
    186.16, 186.1, 186.03, 185.96, 185.9, 185.83, 185.76, 185.69, 185.62, 
    185.56, 185.49, 185.42, 185.35, 185.28, 185.21, 185.14, 185.07, 184.99, 
    184.92, 184.85, 184.78, 184.7, 184.63, 184.55, 184.48, 184.41, 184.33, 
    184.26, 184.18, 184.11, 184.03, 183.96, 183.88, 183.8, 183.73, 183.65, 
    183.58, 183.5, 183.43, 183.36, 183.28, 183.21, 183.13, 183.06, 182.99, 
    182.91, 182.84, 182.77, 182.69, 182.62, 182.55, 182.48, 182.41, 182.34, 
    182.27, 182.2, 182.13, 182.07, 182, 181.94, 181.87, 181.81, 181.75, 
    181.68, 181.62, 181.56, 181.49, 181.43, 181.37, 181.3, 181.24, 181.18, 
    181.12, 181.06, 180.99, 180.93, 180.87, 180.81, 180.75, 180.69, 180.63, 
    180.57, 180.51, 180.45, 180.39, 180.33, 180.27, 180.21, 180.15, 180.09, 
    180.03, 179.97, 179.91, 179.85, 179.79, 179.73, 179.67, 179.6, 179.54, 
    179.47, 179.41, 179.34, 179.28, 179.21, 179.14, 179.08, 179.01, 178.95, 
    178.88, 178.81, 178.75, 178.68, 178.61, 178.55, 178.48, 178.41, 178.35, 
    178.28, 178.22, 178.15, 178.08, 178.01, 177.95, 177.88, 177.81, 177.75, 
    177.68, 177.61, 177.55, 177.48, 177.41, 177.34, 177.27, 177.2, 177.13, 
    177.06, 176.99, 176.92, 176.85, 176.78, 176.72, 176.65, 176.58, 176.51, 
    176.45, 176.38, 176.31, 176.25, 176.18, 176.12, 176.06, 175.99, 175.93, 
    175.86, 175.79, 175.73, 175.66, 175.6, 175.54, 175.47, 175.41, 175.35, 
    175.28, 175.22, 175.16, 175.09, 175.03, 174.97, 174.9, 174.84, 174.78, 
    174.73, 174.67, 174.61, 174.55, 174.49, 174.44, 174.38, 174.32, 174.27, 
    174.21, 174.15, 174.09, 174.03, 173.97, 173.91, 173.85, 173.79, 173.73, 
    173.67, 173.61, 173.55, 173.48, 173.42, 173.36, 173.3, 173.23, 173.17, 
    173.1, 173.04, 172.97, 172.9, 172.84, 172.77, 172.7, 172.64, 172.57, 
    172.5, 172.43, 172.36, 172.29, 172.23, 172.16, 172.09, 172.02, 171.95, 
    171.88, 171.81, 171.75, 171.68, 171.61, 171.54, 171.47, 171.4, 171.33, 
    171.27, 171.2, 171.13, 171.06, 170.99, 170.92, 170.85, 170.78, 170.71, 
    170.64, 170.57, 170.51, 170.44, 170.38, 170.31, 170.24, 170.18, 170.11, 
    170.05, 169.98, 169.91, 169.84, 169.78, 169.71, 169.64, 169.57, 169.5, 
    169.44, 169.37, 169.3, 169.24, 169.17, 169.1, 169.04, 168.97, 168.91, 
    168.84, 168.78, 168.71, 168.65, 168.58, 168.52, 168.45, 168.39, 168.32, 
    168.26, 168.19, 168.13, 168.06, 168, 167.93, 167.87, 167.8, 167.73, 
    167.67, 167.6, 167.53, 167.47, 167.4, 167.33, 167.27, 167.2, 167.14, 
    167.07, 167.01, 166.94, 166.87, 166.81, 166.74, 166.67, 166.61, 166.54, 
    166.47, 166.4, 166.34, 166.27, 166.2, 166.13, 166.06, 165.99, 165.93, 
    165.86, 165.79, 165.72, 165.65, 165.59, 165.52, 165.45, 165.38, 165.31, 
    165.24, 165.17, 165.1, 165.03, 164.97, 164.9, 164.83, 164.77, 164.7, 
    164.64, 164.57, 164.51, 164.44, 164.38, 164.31, 164.25, 164.18, 164.12, 
    164.06, 163.99, 163.93, 163.87, 163.81, 163.75, 163.69, 163.63, 163.57, 
    163.51, 163.45, 163.39, 163.34, 163.28, 163.22, 163.16, 163.11, 163.05, 
    163, 162.94, 162.89, 162.83, 162.77, 162.72, 162.66, 162.61, 162.55, 
    162.49, 162.44, 162.38, 162.32, 162.27, 162.21, 162.15, 162.1, 162.04, 
    161.98, 161.93, 161.87, 161.81, 161.75, 161.7, 161.64, 161.58, 161.52, 
    161.46, 161.41, 161.35, 161.29, 161.23, 161.17, 161.11, 161.05, 160.99, 
    160.93, 160.87, 160.81, 160.75, 160.69, 160.63, 160.57, 160.52, 160.46, 
    160.4, 160.34, 160.28, 160.22, 160.16, 160.11, 160.05, 159.99, 159.93, 
    159.87, 159.81, 159.76, 159.7, 159.64, 159.58, 159.52, 159.47, 159.41, 
    159.35, 159.3, 159.24, 159.18, 159.12, 159.07, 159.01, 158.95, 158.89, 
    158.84, 158.78, 158.72, 158.66, 158.61, 158.55, 158.49, 158.43, 158.37, 
    158.31, 158.25, 158.19, 158.13, 158.07, 158.01, 157.95, 157.89, 157.83, 
    157.77, 157.71, 157.65, 157.59, 157.53, 157.47, 157.41, 157.35, 157.29, 
    157.23, 157.17, 157.1, 157.04, 156.98, 156.92, 156.86, 156.8, 156.74, 
    156.69, 156.63, 156.57, 156.51, 156.46, 156.4, 156.34, 156.28, 156.23, 
    156.17, 156.12, 156.06, 156, 155.95, 155.89, 155.83, 155.78, 155.72, 
    155.66, 155.61, 155.55, 155.49, 155.44, 155.38, 155.33, 155.27, 155.22, 
    155.16, 155.11, 155.05, 155, 154.94, 154.89, 154.83, 154.78, 154.72, 
    154.67, 154.61, 154.56, 154.5, 154.45, 154.39, 154.33, 154.28, 154.22, 
    154.17, 154.11, 154.05, 154, 153.94, 153.89, 153.83, 153.78, 153.72, 
    153.67, 153.61, 153.56, 153.51, 153.45, 153.4, 153.34, 153.29, 153.23, 
    153.18, 153.12, 153.07, 153.01, 152.96, 152.9, 152.85, 152.79, 152.74, 
    152.68, 152.62, 152.57, 152.51, 152.46, 152.4, 152.35, 152.29, 152.23, 
    152.18, 152.12, 152.07, 152.01, 151.96, 151.9, 151.85, 151.79, 151.74, 
    151.68, 151.63, 151.57, 151.52, 151.46, 151.41, 151.35, 151.3, 151.24, 
    151.19, 151.13, 151.08, 151.02, 150.96, 150.91, 150.85, 150.8, 150.74, 
    150.68, 150.62, 150.56, 150.51, 150.45, 150.39, 150.33, 150.27, 150.21, 
    150.15, 150.09, 150.03, 149.97, 149.91, 149.85, 149.79, 149.73, 149.67, 
    149.61, 149.55, 149.49, 149.43, 149.37, 149.31, 149.25, 149.19, 149.13, 
    149.07, 149.01, 148.95, 148.89, 148.83, 148.77, 148.71, 148.65, 148.58, 
    148.52, 148.46, 148.4, 148.34, 148.28, 148.22, 148.16, 148.1, 148.05, 
    147.99, 147.93, 147.87, 147.81, 147.76, 147.7, 147.65, 147.59, 147.53, 
    147.48, 147.42, 147.36, 147.31, 147.25, 147.19, 147.13, 147.08, 147.02, 
    146.97, 146.91, 146.85, 146.8, 146.74, 146.69, 146.63, 146.58, 146.53, 
    146.47, 146.42, 146.37, 146.32, 146.27, 146.21, 146.16, 146.11, 146.06, 
    146.01, 145.95, 145.9, 145.85, 145.79, 145.74, 145.68, 145.63, 145.57, 
    145.52, 145.47, 145.41, 145.36, 145.3, 145.25, 145.19, 145.14, 145.09, 
    145.04, 144.99, 144.93, 144.88, 144.82, 144.77, 144.72, 144.66, 144.61, 
    144.55, 144.5, 144.44, 144.39, 144.33, 144.28, 144.22, 144.16, 144.11, 
    144.05, 144, 143.94, 143.88, 143.83, 143.77, 143.72, 143.66, 143.61, 
    143.55, 143.5, 143.44, 143.39, 143.33, 143.28, 143.22, 143.16, 143.11, 
    143.05, 142.99, 142.93, 142.87, 142.81, 142.76, 142.7, 142.64, 142.58, 
    142.53, 142.47, 142.41, 142.35, 142.29, 142.23, 142.17, 142.11, 142.05, 
    141.99, 141.94, 141.88, 141.82, 141.76, 141.7, 141.64, 141.58, 141.52, 
    141.46, 141.4, 141.34, 141.28, 141.22, 141.16, 141.1, 141.04, 140.98, 
    140.92, 140.86, 140.8, 140.75, 140.69, 140.63, 140.57, 140.51, 140.45, 
    140.39, 140.34, 140.28, 140.22, 140.17, 140.11, 140.06, 140, 139.95, 
    139.9, 139.84, 139.79, 139.74, 139.69, 139.63, 139.58, 139.53, 139.48, 
    139.43, 139.38, 139.33, 139.28, 139.23, 139.18, 139.13, 139.08, 139.03, 
    138.98, 138.93, 138.89, 138.84, 138.79, 138.75, 138.7, 138.66, 138.61, 
    138.57, 138.53, 138.48, 138.44, 138.4, 138.35, 138.31, 138.26, 138.22, 
    138.17, 138.13, 138.09, 138.04, 138, 137.95, 137.91, 137.86, 137.82, 
    137.77, 137.73, 137.68, 137.64, 137.59, 137.54, 137.5, 137.45, 137.41, 
    137.36, 137.32, 137.27, 137.22, 137.18, 137.13, 137.08, 137.03, 136.99, 
    136.94, 136.89, 136.84, 136.79, 136.74, 136.69, 136.64, 136.59, 136.54, 
    136.49, 136.44, 136.39, 136.34, 136.29, 136.24, 136.19, 136.14, 136.09, 
    136.04, 135.99, 135.94, 135.88, 135.83, 135.78, 135.73, 135.68, 135.63, 
    135.58, 135.52, 135.47, 135.42, 135.37, 135.31, 135.26, 135.21, 135.15, 
    135.1, 135.05, 134.99, 134.94, 134.89, 134.83, 134.78, 134.73, 134.68, 
    134.62, 134.57, 134.52, 134.46, 134.41, 134.35, 134.3, 134.24, 134.19, 
    134.13, 134.07, 134.02, 133.96, 133.91, 133.85, 133.8, 133.75, 133.69, 
    133.64, 133.58, 133.53, 133.47, 133.42, 133.37, 133.31, 133.26, 133.2, 
    133.15, 133.09, 133.04, 132.98, 132.93, 132.88, 132.82, 132.76, 132.71, 
    132.65, 132.6, 132.54, 132.49, 132.43, 132.38, 132.32, 132.27, 132.21, 
    132.16, 132.11, 132.06, 132, 131.95, 131.9, 131.85, 131.8, 131.74, 
    131.69, 131.64, 131.58, 131.53, 131.48, 131.42, 131.37, 131.32, 131.27, 
    131.21, 131.16, 131.11, 131.05, 131, 130.95, 130.9, 130.84, 130.79, 
    130.74, 130.69, 130.64, 130.59, 130.54, 130.48, 130.43, 130.38, 130.33, 
    130.28, 130.23, 130.18, 130.13, 130.08, 130.02, 129.97, 129.92, 129.86, 
    129.81, 129.76, 129.7, 129.65, 129.6, 129.54, 129.49, 129.43, 129.38, 
    129.32, 129.27, 129.22, 129.17, 129.12, 129.06, 129.01, 128.96, 128.91, 
    128.86, 128.8, 128.75, 128.7, 128.65, 128.6, 128.55, 128.49, 128.44, 
    128.39, 128.33, 128.28, 128.23, 128.17, 128.12, 128.07, 128.02, 127.97, 
    127.92, 127.86, 127.81, 127.76, 127.71, 127.66, 127.61, 127.56, 127.51, 
    127.46, 127.42, 127.37, 127.32, 127.27, 127.22, 127.17, 127.12, 127.07, 
    127.02, 126.97, 126.92, 126.87, 126.82, 126.77, 126.72, 126.67, 126.62, 
    126.57, 126.53, 126.48, 126.43, 126.38, 126.33, 126.29, 126.24, 126.19, 
    126.14, 126.09, 126.04, 125.99, 125.94, 125.89, 125.84, 125.79, 125.74, 
    125.69, 125.65, 125.6, 125.55, 125.5, 125.45, 125.4, 125.36, 125.31, 
    125.26, 125.21, 125.17, 125.12, 125.07, 125.02, 124.98, 124.93, 124.88, 
    124.83, 124.79, 124.74, 124.69, 124.64, 124.59, 124.53, 124.48, 124.43, 
    124.38, 124.33, 124.28, 124.23, 124.18, 124.13, 124.08, 124.03, 123.98, 
    123.93, 123.88, 123.83, 123.78, 123.73, 123.68, 123.63, 123.58, 123.53, 
    123.48, 123.43, 123.38, 123.33, 123.28, 123.23, 123.18, 123.13, 123.08, 
    123.03, 122.98, 122.93, 122.88, 122.83, 122.78, 122.73, 122.68, 122.63, 
    122.58, 122.53, 122.48, 122.43, 122.39, 122.34, 122.29, 122.25, 122.2, 
    122.15, 122.1, 122.05, 122.01, 121.96, 121.91, 121.86, 121.82, 121.77, 
    121.72, 121.67, 121.63, 121.58, 121.53, 121.48, 121.43, 121.39, 121.34, 
    121.29, 121.24, 121.2, 121.15, 121.1, 121.05, 121.01, 120.96, 120.91, 
    120.87, 120.83, 120.78, 120.74, 120.69, 120.65, 120.6, 120.56, 120.51, 
    120.46, 120.42, 120.37, 120.33, 120.28, 120.23, 120.19, 120.14, 120.09, 
    120.05, 120, 119.96, 119.91, 119.87, 119.82, 119.78, 119.73, 119.69, 
    119.65, 119.6, 119.56, 119.52, 119.48, 119.43, 119.39, 119.35, 119.3, 
    119.26, 119.21, 119.17, 119.13, 119.08, 119.04, 119, 118.95, 118.91, 
    118.86, 118.82, 118.78, 118.73, 118.69, 118.64, 118.6, 118.55, 118.51, 
    118.47, 118.42, 118.38, 118.34, 118.29, 118.24, 118.2, 118.15, 118.1, 
    118.06, 118.01, 117.96, 117.91, 117.86, 117.82, 117.77, 117.72, 117.67, 
    117.63, 117.58, 117.53, 117.49, 117.44, 117.4, 117.35, 117.31, 117.26, 
    117.22, 117.17, 117.12, 117.08, 117.03, 116.99, 116.94, 116.9, 116.85, 
    116.81, 116.77, 116.72, 116.68, 116.63, 116.59, 116.55, 116.5, 116.46, 
    116.42, 116.37, 116.33, 116.29, 116.25, 116.21, 116.16, 116.12, 116.08, 
    116.04, 116, 115.96, 115.92, 115.88, 115.84, 115.8, 115.76, 115.71, 
    115.67, 115.63, 115.59, 115.54, 115.5, 115.46, 115.41, 115.37, 115.33, 
    115.28, 115.24, 115.19, 115.15, 115.1, 115.06, 115.01, 114.97, 114.93, 
    114.88, 114.84, 114.79, 114.75, 114.7, 114.66, 114.61, 114.57, 114.52, 
    114.47, 114.43, 114.38, 114.34, 114.29, 114.24, 114.2, 114.15, 114.1, 
    114.05, 114.01, 113.96, 113.91, 113.87, 113.82, 113.77, 113.72, 113.68, 
    113.63, 113.58, 113.53, 113.49, 113.44, 113.39, 113.35, 113.3, 113.25, 
    113.21, 113.16, 113.12, 113.07, 113.03, 112.98, 112.94, 112.89, 112.85, 
    112.81, 112.76, 112.72, 112.67, 112.63, 112.58, 112.54, 112.49, 112.45, 
    112.4, 112.36, 112.32, 112.27, 112.23, 112.18, 112.14, 112.09, 112.05, 
    112, 111.96, 111.92, 111.87, 111.83, 111.79, 111.75, 111.71, 111.66, 
    111.62, 111.58, 111.54, 111.49, 111.45, 111.41, 111.36, 111.32, 111.27, 
    111.23, 111.19, 111.14, 111.1, 111.06, 111.01, 110.97, 110.93, 110.89, 
    110.85, 110.81, 110.77, 110.72, 110.68, 110.64, 110.6, 110.55, 110.51, 
    110.47, 110.43, 110.39, 110.34, 110.3, 110.26, 110.22, 110.17, 110.13, 
    110.09, 110.04, 110, 109.95, 109.91, 109.86, 109.82, 109.77, 109.73, 
    109.68, 109.63, 109.59, 109.54, 109.5, 109.45, 109.41, 109.36, 109.32, 
    109.27, 109.23, 109.18, 109.13, 109.09, 109.04, 108.99, 108.95, 108.9, 
    108.85, 108.81, 108.76, 108.71, 108.66, 108.61, 108.57, 108.52, 108.47, 
    108.42, 108.38, 108.33, 108.28, 108.24, 108.19, 108.15, 108.1, 108.06, 
    108.01, 107.97, 107.92, 107.88, 107.83, 107.79, 107.74, 107.69, 107.65, 
    107.6, 107.55, 107.51, 107.46, 107.41, 107.37, 107.32, 107.28, 107.23, 
    107.19, 107.14, 107.1, 107.06, 107.02, 106.97, 106.93, 106.89, 106.85, 
    106.81, 106.77, 106.73, 106.69, 106.65, 106.61, 106.57, 106.53, 106.48, 
    106.44, 106.4, 106.36, 106.32, 106.28, 106.24, 106.2, 106.16, 106.12, 
    106.08, 106.04, 106, 105.96, 105.92, 105.89, 105.85, 105.81, 105.77, 
    105.73, 105.69, 105.65, 105.61, 105.57, 105.53, 105.49, 105.45, 105.41, 
    105.37, 105.33, 105.29, 105.25, 105.21, 105.17, 105.14, 105.1, 105.06, 
    105.02, 104.98, 104.95, 104.91, 104.87, 104.83, 104.79, 104.76, 104.72, 
    104.68, 104.64, 104.6, 104.56, 104.52, 104.49, 104.45, 104.41, 104.37, 
    104.33, 104.29, 104.26, 104.22, 104.18, 104.14, 104.1, 104.06, 104.02, 
    103.98, 103.95, 103.91, 103.87, 103.83, 103.79, 103.75, 103.71, 103.67, 
    103.63, 103.59, 103.55, 103.51, 103.47, 103.43, 103.39, 103.35, 103.31, 
    103.27, 103.23, 103.19, 103.15, 103.11, 103.07, 103.03, 102.99, 102.95, 
    102.9, 102.86, 102.82, 102.78, 102.74, 102.7, 102.66, 102.62, 102.58, 
    102.54, 102.5, 102.46, 102.42, 102.37, 102.33, 102.29, 102.25, 102.21, 
    102.17, 102.13, 102.08, 102.04, 102, 101.95, 101.91, 101.87, 101.83, 
    101.78, 101.74, 101.7, 101.66, 101.61, 101.57, 101.52, 101.48, 101.44, 
    101.39, 101.35, 101.31, 101.26, 101.22, 101.18, 101.14, 101.09, 101.05, 
    101.01, 100.97, 100.93, 100.88, 100.84, 100.8, 100.76, 100.72, 100.68, 
    100.64, 100.59, 100.55, 100.51, 100.47, 100.43, 100.39, 100.35, 100.31, 
    100.27, 100.22, 100.18, 100.14, 100.1, 100.06, 100.02, 99.98, 99.939, 
    99.898, 99.858, 99.817, 99.776, 99.734, 99.693, 99.652, 99.61, 99.569, 
    99.527, 99.485, 99.443, 99.4, 99.358, 99.315, 99.273, 99.231, 99.189, 
    99.146, 99.104, 99.062, 99.019, 98.977, 98.935, 98.894, 98.852, 98.81, 
    98.768, 98.726, 98.684, 98.642, 98.6, 98.558, 98.517, 98.475, 98.433, 
    98.391, 98.349, 98.306, 98.264, 98.221, 98.179, 98.137, 98.094, 98.052, 
    98.01, 97.967, 97.925, 97.883, 97.842, 97.8, 97.758, 97.715, 97.673, 
    97.629, 97.586, 97.543, 97.5, 97.457, 97.414, 97.37, 97.327, 97.283, 
    97.24, 97.197, 97.154, 97.111, 97.068, 97.026, 96.984, 96.943, 96.902, 
    96.861, 96.82, 96.78, 96.74, 96.701, 96.662, 96.622, 96.583, 96.544, 
    96.504, 96.464, 96.424, 96.383, 96.342, 96.301, 96.26, 96.22, 96.179, 
    96.139, 96.098, 96.058, 96.018, 95.977, 95.938, 95.898, 95.859, 95.821, 
    95.782, 95.744, 95.705, 95.667, 95.629, 95.59, 95.552, 95.514, 95.476, 
    95.438, 95.399, 95.36, 95.321, 95.282, 95.242, 95.203, 95.163, 95.124, 
    95.084, 95.045, 95.006, 94.968, 94.93, 94.892, 94.855, 94.818, 94.78, 
    94.742, 94.704, 94.667, 94.629, 94.591, 94.553, 94.515, 94.477, 94.438, 
    94.4, 94.362, 94.324, 94.286, 94.249, 94.212, 94.175, 94.138, 94.101, 
    94.063, 94.025, 93.986, 93.947, 93.909, 93.87, 93.831, 93.792, 93.753, 
    93.713, 93.674, 93.634, 93.595, 93.557, 93.518, 93.479, 93.44, 93.402, 
    93.363, 93.325, 93.286, 93.248, 93.21, 93.173, 93.135, 93.097, 93.06, 
    93.022, 92.984, 92.946, 92.907, 92.868, 92.829, 92.789, 92.749, 92.708, 
    92.667, 92.626, 92.586, 92.545, 92.505, 92.466, 92.427, 92.388, 92.349, 
    92.311, 92.272, 92.234, 92.196, 92.158, 92.12, 92.082, 92.044, 92.006, 
    91.969, 91.931, 91.894, 91.857, 91.818, 91.78, 91.741, 91.702, 91.664, 
    91.626, 91.588, 91.55, 91.512, 91.475, 91.437, 91.399, 91.362, 91.324, 
    91.287, 91.251, 91.214, 91.177, 91.14, 91.103, 91.066, 91.029, 90.992, 
    90.955, 90.918, 90.881, 90.843, 90.804, 90.766, 90.728, 90.689, 90.651, 
    90.613, 90.574, 90.535, 90.495, 90.455, 90.416, 90.378, 90.34, 90.302, 
    90.264, 90.226, 90.188, 90.15, 90.111, 90.072, 90.033, 89.995, 89.957, 
    89.919, 89.881, 89.843, 89.805, 89.768, 89.731, 89.695, 89.658, 89.622, 
    89.586, 89.55, 89.514, 89.479, 89.444, 89.409, 89.374, 89.339, 89.304, 
    89.269, 89.234, 89.199, 89.165, 89.13, 89.095, 89.06, 89.026, 88.991, 
    88.957, 88.922, 88.888, 88.854, 88.82, 88.786, 88.753, 88.719, 88.685, 
    88.651, 88.617, 88.582, 88.546, 88.51, 88.474, 88.437, 88.4, 88.362, 
    88.325, 88.288, 88.25, 88.213, 88.176, 88.138, 88.1, 88.063, 88.025, 
    87.987, 87.95, 87.912, 87.874, 87.836, 87.798, 87.759, 87.72, 87.681, 
    87.642, 87.602, 87.562, 87.522, 87.482, 87.441, 87.4, 87.358, 87.316, 
    87.274, 87.232, 87.19, 87.148, 87.106, 87.064, 87.023, 86.981, 86.94, 
    86.898, 86.855, 86.813, 86.77, 86.727, 86.685, 86.642, 86.599, 86.556, 
    86.514, 86.471, 86.427, 86.384, 86.34, 86.296, 86.251, 86.207, 86.161, 
    86.116, 86.07, 86.025, 85.979, 85.933, 85.888, 85.842, 85.796, 85.751, 
    85.706, 85.662, 85.618, 85.574, 85.53, 85.486, 85.441, 85.396, 85.351, 
    85.305, 85.26, 85.215, 85.17, 85.124, 85.078, 85.032, 84.985, 84.938, 
    84.891, 84.844, 84.796, 84.749, 84.702, 84.655, 84.608, 84.562, 84.517, 
    84.472, 84.427, 84.382, 84.338, 84.293, 84.249, 84.204, 84.159, 84.113, 
    84.067, 84.021, 83.973, 83.926, 83.878, 83.83, 83.782, 83.734, 83.686, 
    83.638, 83.59, 83.543, 83.495, 83.447, 83.399, 83.351, 83.303, 83.254, 
    83.206, 83.157, 83.109, 83.06, 83.011, 82.962, 82.912, 82.862, 82.812, 
    82.762, 82.712, 82.662, 82.611, 82.561, 82.51, 82.459, 82.409, 82.358, 
    82.307, 82.257, 82.206, 82.156, 82.105, 82.054, 82.003, 81.952, 81.901, 
    81.849, 81.797, 81.746, 81.695, 81.644, 81.593, 81.542, 81.492, 81.442, 
    81.392, 81.342, 81.292, 81.242, 81.192, 81.142, 81.091, 81.039, 80.987, 
    80.935, 80.883, 80.83, 80.777, 80.724, 80.67, 80.616, 80.562, 80.508, 
    80.454, 80.4, 80.346, 80.292, 80.238, 80.184, 80.131, 80.079, 80.027, 
    79.976, 79.925, 79.876, 79.827, 79.778, 79.729, 79.68, 79.632, 79.584, 
    79.537, 79.489, 79.442, 79.396, 79.35, 79.304, 79.26, 79.216, 79.173, 
    79.132, 79.091, 79.051, 79.011, 78.972, 78.933, 78.896, 78.858, 78.822, 
    78.785, 78.748, 78.712, 78.676, 78.641, 78.607, 78.573, 78.539, 78.505, 
    78.471, 78.436, 78.402, 78.368, 78.334, 78.3, 78.266, 78.231, 78.197, 
    78.162, 78.128, 78.093, 78.058, 78.022, 77.987, 77.951, 77.914, 77.878, 
    77.84, 77.803, 77.766, 77.729, 77.691, 77.654, 77.617, 77.581, 77.544, 
    77.508, 77.473, 77.438, 77.404, 77.369, 77.334, 77.299, 77.265, 77.23, 
    77.195, 77.161, 77.126, 77.092, 77.058, 77.024, 76.989, 76.954, 76.918, 
    76.883, 76.849, 76.815, 76.781, 76.747, 76.713, 76.679, 76.645, 76.612, 
    76.578, 76.546, 76.513, 76.48, 76.447, 76.414, 76.381, 76.348, 76.314, 
    76.28, 76.246, 76.211, 76.176, 76.141, 76.105, 76.07, 76.033, 75.997, 
    75.96, 75.922, 75.884, 75.846, 75.807, 75.767, 75.726, 75.685, 75.644, 
    75.602, 75.56, 75.518, 75.474, 75.43, 75.385, 75.34, 75.295, 75.25, 
    75.206, 75.161, 75.116, 75.071, 75.027, 74.982, 74.938, 74.893, 74.849, 
    74.805, 74.76, 74.715, 74.671, 74.626, 74.581, 74.536, 74.491, 74.446, 
    74.401, 74.355, 74.311, 74.266, 74.222, 74.178, 74.135, 74.092, 74.048, 
    74.005, 73.963, 73.92, 73.878, 73.836, 73.795, 73.753, 73.711, 73.67, 
    73.628, 73.587, 73.545, 73.503, 73.461, 73.418, 73.376, 73.333, 73.289, 
    73.245, 73.201, 73.156, 73.111, 73.066, 73.019, 72.972, 72.924, 72.877, 
    72.829, 72.782, 72.734, 72.687, 72.64, 72.593, 72.547, 72.5, 72.455, 
    72.409, 72.365, 72.321, 72.278, 72.235, 72.192, 72.149, 72.106, 72.063, 
    72.019, 71.976, 71.933, 71.89, 71.847, 71.804, 71.762, 71.719, 71.677, 
    71.635, 71.594, 71.553, 71.513, 71.474, 71.435, 71.398, 71.36, 71.323, 
    71.286, 71.25, 71.212, 71.175, 71.137, 71.098, 71.058, 71.018, 70.976, 
    70.935, 70.892, 70.849, 70.806, 70.762, 70.718, 70.673, 70.628, 70.583, 
    70.539, 70.494, 70.45, 70.406, 70.361, 70.316, 70.272, 70.227, 70.181, 
    70.136, 70.091, 70.046, 70, 69.954, 69.908, 69.862, 69.815, 69.769, 
    69.723, 69.678, 69.633, 69.589, 69.545, 69.502, 69.459, 69.416, 69.373, 
    69.331, 69.289, 69.247, 69.205, 69.162, 69.119, 69.076, 69.033, 68.99, 
    68.947, 68.905, 68.862, 68.819, 68.777, 68.734, 68.691, 68.648, 68.606, 
    68.563, 68.52, 68.477, 68.434, 68.39, 68.346, 68.302, 68.258, 68.214, 
    68.169, 68.124, 68.079, 68.034, 67.988, 67.942, 67.895, 67.849, 67.803, 
    67.757, 67.711, 67.667, 67.623, 67.581, 67.539, 67.497, 67.456, 67.416, 
    67.376, 67.335, 67.295, 67.255, 67.214, 67.174, 67.133, 67.093, 67.052, 
    67.011, 66.97, 66.929, 66.888, 66.847, 66.806, 66.765, 66.725, 66.684, 
    66.644, 66.603, 66.563, 66.522, 66.481, 66.44, 66.4, 66.359, 66.32, 
    66.28, 66.241, 66.202, 66.162, 66.123, 66.084, 66.045, 66.006, 65.967, 
    65.928, 65.89, 65.851, 65.813, 65.775, 65.738, 65.7, 65.663, 65.626, 
    65.59, 65.554, 65.519, 65.483, 65.448, 65.413, 65.378, 65.344, 65.31, 
    65.276, 65.243, 65.21, 65.178, 65.147, 65.116, 65.085, 65.054, 65.023, 
    64.993, 64.962, 64.932, 64.901, 64.87, 64.839, 64.807, 64.775, 64.742, 
    64.709, 64.675, 64.641, 64.607, 64.572, 64.537, 64.502, 64.466, 64.429, 
    64.392, 64.354, 64.317, 64.279, 64.242, 64.205, 64.168, 64.131, 64.094, 
    64.057, 64.021, 63.984, 63.947, 63.91, 63.873, 63.835, 63.798, 63.76, 
    63.722, 63.684, 63.646, 63.607, 63.569, 63.53, 63.491, 63.451, 63.412, 
    63.373, 63.335, 63.297, 63.259, 63.22, 63.182, 63.144, 63.106, 63.068, 
    63.031, 62.994, 62.958, 62.922, 62.886, 62.85, 62.814, 62.777, 62.741, 
    62.704, 62.667, 62.63, 62.592, 62.554, 62.516, 62.478, 62.439, 62.4, 
    62.362, 62.323, 62.283, 62.244, 62.205, 62.166, 62.127, 62.089, 62.051, 
    62.013, 61.975, 61.937, 61.899, 61.862, 61.824, 61.787, 61.749, 61.712, 
    61.675, 61.639, 61.603, 61.567, 61.531, 61.495, 61.46, 61.426, 61.392, 
    61.358, 61.325, 61.293, 61.26, 61.228, 61.195, 61.163, 61.131, 61.098, 
    61.066, 61.034, 61.002, 60.969, 60.937, 60.905, 60.872, 60.839, 60.807, 
    60.774, 60.741, 60.708, 60.676, 60.643, 60.61, 60.578, 60.545, 60.513, 
    60.481, 60.448, 60.416, 60.383, 60.351, 60.318, 60.286, 60.253, 60.22, 
    60.186, 60.153, 60.118, 60.084, 60.049, 60.014, 59.979, 59.943, 59.908, 
    59.873, 59.837, 59.802, 59.767, 59.733, 59.698, 59.664, 59.63, 59.597, 
    59.563, 59.53, 59.496, 59.463, 59.429, 59.395, 59.36, 59.325, 59.29, 
    59.255, 59.22, 59.185, 59.15, 59.115, 59.08, 59.045, 59.01, 58.976, 
    58.942, 58.907, 58.873, 58.839, 58.806, 58.772, 58.739, 58.705, 58.672, 
    58.639, 58.606, 58.573, 58.54, 58.507, 58.474, 58.442, 58.41, 58.378, 
    58.346, 58.314, 58.282, 58.251, 58.219, 58.188, 58.157, 58.127, 58.097, 
    58.067, 58.037, 58.008, 57.978, 57.949, 57.92, 57.891, 57.862, 57.833, 
    57.804, 57.775, 57.745, 57.716, 57.686, 57.656, 57.626, 57.596, 57.566, 
    57.537, 57.507, 57.478, 57.449, 57.421, 57.393, 57.366, 57.34, 57.315, 
    57.211, 57.109, 57.01, 56.912, 56.816, 56.722, 56.629, 56.537, 56.447, 
    56.356, 56.266, 56.175, 56.084, 55.992, 55.899, 55.804, 55.708, 55.61, 
    55.51, 55.407, 55.303, 55.197, 55.089, 54.979, 54.868, 54.755, 54.641, 
    54.527, 54.411, 54.296, 54.181, 54.066, 53.952, 53.839, 53.726, 53.615, 
    53.505, 53.397, 53.29, 53.184, 53.08, 52.977, 52.875, 52.774, 52.674, 
    52.574, 52.475, 52.376, 52.277, 52.179, 52.08, 51.98, 51.88, 51.78, 
    51.679, 51.578, 51.476, 51.373, 51.269, 51.165, 51.061, 50.955, 50.85, 
    50.744, 50.638, 50.532, 50.426, 50.32, 50.215, 50.11, 50.005, 49.901, 
    49.798, 49.695, 49.593, 49.491, 49.39, 49.29, 49.19, 49.09, 48.991, 
    48.892, 48.793, 48.694, 48.595, 48.496, 48.396, 48.296, 48.195, 48.095, 
    47.993, 47.892, 47.789, 47.687, 47.584, 47.481, 47.377, 47.274, 47.17, 
    47.066, 46.962, 46.858, 46.754, 46.65, 46.547, 46.443, 46.34, 46.236, 
    46.133, 46.03, 45.928, 45.825, 45.723, 45.621, 45.52, 45.419, 45.318, 
    45.218, 45.118, 45.018, 44.919, 44.821, 44.723, 44.625, 44.528, 44.432, 
    44.336, 44.24, 44.145, 44.051, 43.957, 43.863, 43.77, 43.677, 43.585, 
    43.493, 43.401, 43.309, 43.218, 43.126, 43.035, 42.944, 42.852, 42.761, 
    42.669, 42.577, 42.484, 42.392, 42.298, 42.204, 42.11, 42.015, 41.92, 
    41.824, 41.728, 41.631, 41.533, 41.436, 41.338, 41.24, 41.141, 41.042, 
    40.944, 40.845, 40.746, 40.647, 40.548, 40.449, 40.351, 40.252, 40.154, 
    40.056, 39.958, 39.86, 39.763, 39.666, 39.57, 39.473, 39.377, 39.281, 
    39.186, 39.091, 38.996, 38.901, 38.807, 38.713, 38.619, 38.526, 38.432, 
    38.339, 38.247, 38.154, 38.062, 37.97, 37.878, 37.786, 37.695, 37.604, 
    37.513, 37.422, 37.331, 37.24, 37.149, 37.057, 36.966, 36.873, 36.781, 
    36.688, 36.594, 36.499, 36.403, 36.307, 36.209, 36.11, 36.011, 35.91, 
    35.808, 35.705, 35.601, 35.497, 35.391, 35.285, 35.178, 35.07, 34.962, 
    34.854, 34.745, 34.636, 34.527, 34.418, 34.309, 34.2, 34.092, 33.983, 
    33.874, 33.766, 33.658, 33.55, 33.442, 33.335, 33.228, 33.12, 33.014, 
    32.907, 32.8, 32.694, 32.588, 32.482, 32.377, 32.272, 32.168, 32.064, 
    31.961, 31.859, 31.757, 31.657, 31.557, 31.459, 31.362, 31.266, 31.171, 
    31.078, 30.986, 30.895, 30.806, 30.718, 30.631, 30.545, 30.461, 30.378, 
    30.296, 30.215, 30.135, 30.056, 29.977, 29.899, 29.821, 29.744, 29.667, 
    29.59, 29.514, 29.437, 29.361, 29.285, 29.209, 29.133, 29.057, 28.982, 
    28.906, 28.831, 28.756, 28.681, 28.607, 28.533, 28.459, 28.385, 28.312, 
    28.239, 28.165, 28.092, 28.019, 27.946, 27.873, 27.799, 27.725, 27.651, 
    27.576, 27.501, 27.425, 27.349, 27.273, 27.195, 27.117, 27.039, 26.96, 
    26.88, 26.8, 26.719, 26.638, 26.556, 26.473, 26.39, 26.306, 26.222, 
    26.137, 26.052, 25.967, 25.88, 25.794, 25.707, 25.62, 25.532, 25.444, 
    25.355, 25.267, 25.178, 25.089, 25, 24.91, 24.821, 24.731, 24.642, 
    24.553, 24.463, 24.374, 24.285, 24.197, 24.108, 24.02, 23.932, 23.844, 
    23.757, 23.67, 23.583, 23.497, 23.411, 23.326, 23.241, 23.157, 23.073, 
    22.99, 22.907, 22.825, 22.743, 22.661, 22.58, 22.5, 22.42, 22.341, 
    22.262, 22.184, 22.106, 22.028, 21.951, 21.874, 21.798, 21.723, 21.647, 
    21.572, 21.497, 21.423, 21.349, 21.276, 21.202, 21.13, 21.057, 20.985, 
    20.913, 20.841, 20.77, 20.699, 20.629, 20.559, 20.489, 20.42, 20.35, 
    20.282, 20.213, 20.145, 20.076, 20.008, 19.94, 19.872, 19.804, 19.736, 
    19.668, 19.599, 19.531, 19.462, 19.393, 19.324, 19.254, 19.184, 19.114, 
    19.044, 18.974, 18.904, 18.833, 18.763, 18.693, 18.622, 18.552, 18.482, 
    18.413, 18.343, 18.274, 18.205, 18.137, 18.069, 18.001, 17.934, 17.867, 
    17.8, 17.734, 17.668, 17.602, 17.536, 17.471, 17.406, 17.342, 17.277, 
    17.213, 17.148, 17.084, 17.02, 16.956, 16.892, 16.829, 16.765, 16.702, 
    16.638, 16.575, 16.512, 16.45, 16.387, 16.324, 16.262, 16.2, 16.138, 
    16.076, 16.014, 15.952, 15.89, 15.828, 15.766, 15.704, 15.642, 15.579, 
    15.516, 15.454, 15.39, 15.327, 15.264, 15.2, 15.136, 15.072, 15.008, 
    14.943, 14.879, 14.814, 14.75, 14.685, 14.621, 14.556, 14.492, 14.428, 
    14.364, 14.301, 14.238, 14.175, 14.112, 14.05, 13.988, 13.927, 13.866, 
    13.806, 13.746, 13.687, 13.629, 13.571, 13.514, 13.457, 13.401, 13.346, 
    13.291, 13.237, 13.183, 13.13, 13.078, 13.026, 12.974, 12.923, 12.872, 
    12.821, 12.77, 12.72, 12.669, 12.619, 12.569, 12.519, 12.468, 12.418, 
    12.367, 12.317, 12.266, 12.215, 12.164, 12.112, 12.061, 12.009, 11.957, 
    11.905, 11.853, 11.801, 11.748, 11.696, 11.643, 11.591, 11.538, 11.486, 
    11.433, 11.381, 11.329, 11.277, 11.225, 11.173, 11.121, 11.07, 11.018, 
    10.967, 10.916, 10.865, 10.814, 10.763, 10.713, 10.662, 10.612, 10.562, 
    10.512, 10.462, 10.412, 10.362, 10.313, 10.263, 10.214, 10.165, 10.116, 
    10.067, 10.019, 9.9709, 9.9232, 9.8759, 9.8289, 9.7823, 9.7361, 9.6903, 
    9.6449, 9.6, 9.5554, 9.5112, 9.4674, 9.4239, 9.3807, 9.3379, 9.2954, 
    9.2531, 9.2111, 9.1693, 9.1277, 9.0863, 9.045, 9.0039, 8.963, 8.9222, 
    8.8815, 8.8409, 8.8004, 8.76, 8.7197, 8.6794, 8.6393, 8.5991, 8.5591, 
    8.519, 8.479, 8.439, 8.399, 8.359, 8.3191, 8.2791, 8.2391, 8.1991, 
    8.1591, 8.1191, 8.0791, 8.0391, 7.9991, 7.9592, 7.9193, 7.8795, 7.8398, 
    7.8002, 7.7606, 7.7211, 7.6818, 7.6426, 7.6035, 7.5645, 7.5256, 7.4868, 
    7.4482, 7.4097, 7.3713, 7.3331, 7.2949, 7.2569, 7.219, 7.1813, 7.1437, 
    7.1063, 7.069, 7.0318, 6.9948, 6.958, 6.9214, 6.8849, 6.8486, 6.8124, 
    6.7765, 6.7406, 6.705, 6.6695, 6.6341, 6.5988, 6.5637, 6.5287, 6.4939, 
    6.4592, 6.4246, 6.3902, 6.3559, 6.3218, 6.2879, 6.2542, 6.2208, 6.1876, 
    6.1546, 6.1219, 6.0896, 6.0575, 6.0257, 5.9943, 5.9631, 5.9323, 5.9018, 
    5.8715, 5.8416, 5.8119, 5.7825, 5.7534, 5.7245, 5.6958, 5.6674, 5.6392, 
    5.6111, 5.5832, 5.5556, 5.528, 5.5006, 5.4734, 5.4463, 5.4192, 5.3923, 
    5.3655, 5.3387, 5.312, 5.2853, 5.2587, 5.232, 5.2054, 5.1787, 5.1521, 
    5.1254, 5.0986, 5.0718, 5.045, 5.0181, 4.9912, 4.9643, 4.9372, 4.9102, 
    4.8831, 4.856, 4.8289, 4.8018, 4.7748, 4.7477, 4.7207, 4.6937, 4.6667, 
    4.6398, 4.613, 4.5863, 4.5596, 4.5331, 4.5066, 4.4802, 4.454, 4.4278, 
    4.4018, 4.3759, 4.3501, 4.3244, 4.2988, 4.2734, 4.2481, 4.2229, 4.1979, 
    4.173, 4.1482, 4.1235, 4.099, 4.0746, 4.0503, 4.0262, 4.0022, 3.9783, 
    3.9546, 3.9309, 3.9074, 3.8841, 3.8608, 3.8377, 3.8147, 3.7918, 3.7691, 
    3.7464, 3.7239, 3.7016, 3.6793, 3.6572, 3.6353, 3.6134, 3.5917, 3.5701, 
    3.5487, 3.5274, 3.5062, 3.4852, 3.4644, 3.4437, 3.4232, 3.4028, 3.3826, 
    3.3626, 3.3428, 3.3232, 3.3037, 3.2845, 3.2654, 3.2465, 3.2279, 3.2094, 
    3.191, 3.1729, 3.1549, 3.1371, 3.1195, 3.102, 3.0846, 3.0674, 3.0503, 
    3.0333, 3.0164, 2.9997, 2.983, 2.9664, 2.9499, 2.9334, 2.917, 2.9006, 
    2.8843, 2.8681, 2.8518, 2.8357, 2.8195, 2.8034, 2.7873, 2.7713, 2.7553, 
    2.7393, 2.7234, 2.7075, 2.6917, 2.6759, 2.6602, 2.6446, 2.6291, 2.6136, 
    2.5982, 2.5829, 2.5676, 2.5525, 2.5375, 2.5226, 2.5077, 2.493, 2.4784, 
    2.4639, 2.4496, 2.4353, 2.4212, 2.4072, 2.3933, 2.3795, 2.3658, 2.3522, 
    2.3388, 2.3254, 2.3121, 2.2989, 2.2859, 2.2729, 2.2599, 2.2471, 2.2343, 
    2.2216, 2.2089, 2.1964, 2.1838, 2.1714, 2.159, 2.1466, 2.1343, 2.1221, 
    2.11, 2.0979, 2.0859, 2.0739, 2.062, 2.0502, 2.0385, 2.0268, 2.0152, 
    2.0037, 1.9922, 1.9808, 1.9695, 1.9582, 1.947, 1.9359, 1.9248, 1.9137, 
    1.9027, 1.8918, 1.8809, 1.8701, 1.8592, 1.8484, 1.8377, 1.8269, 1.8162, 
    1.8056, 1.7949, 1.7842, 1.7736, 1.763, 1.7524, 1.7419, 1.7313, 1.7208, 
    1.7103, 1.6998, 1.6894, 1.679, 1.6686, 1.6583, 1.648, 1.6378, 1.6276, 
    1.6175, 1.6074, 1.5974, 1.5874, 1.5775, 1.5677, 1.5579, 1.5482, 1.5386, 
    1.529, 1.5195, 1.5101, 1.5007, 1.4914, 1.4822, 1.4731, 1.4641, 1.4551, 
    1.4462, 1.4374, 1.4286, 1.42, 1.4114, 1.4029, 1.3945, 1.3861, 1.3778, 
    1.3696, 1.3615, 1.3534, 1.3454, 1.3374, 1.3296, 1.3217, 1.3139, 1.3062, 
    1.2985, 1.2908, 1.2832, 1.2756, 1.268, 1.2605, 1.253, 1.2456, 1.2382, 
    1.2308, 1.2235, 1.2162, 1.209, 1.2018, 1.1947, 1.1877, 1.1807, 1.1738, 
    1.1669, 1.1601, 1.1534, 1.1467, 1.1401, 1.1336, 1.1271, 1.1207, 1.1143, 
    1.108, 1.1017, 1.0955, 1.0893, 1.0831, 1.077, 1.0708, 1.0647, 1.0586, 
    1.0526, 1.0465, 1.0405, 1.0345, 1.0284, 1.0224, 1.0164, 1.0104, 1.0044, 
    0.99844, 0.99248, 0.98652, 0.98057, 0.97464, 0.96873, 0.96284, 0.95697, 
    0.95112, 0.9453, 0.93951, 0.93376, 0.92803, 0.92235, 0.9167, 0.9111, 
    0.90554, 0.90003, 0.89457, 0.88916, 0.88381, 0.87851, 0.87326, 0.86806, 
    0.86293, 0.85785, 0.85282, 0.84786, 0.84294, 0.83809, 0.83328, 0.82853, 
    0.82383, 0.81918, 0.81458, 0.81002, 0.80551, 0.80104, 0.7966, 0.79221, 
    0.78785, 0.78352, 0.77922, 0.77495, 0.7707, 0.76648, 0.76227, 0.75809, 
    0.75392, 0.74976, 0.74562, 0.74148, 0.73736, 0.73325, 0.72915, 0.72505, 
    0.72097, 0.71689, 0.71283, 0.70877, 0.70473, 0.7007, 0.69668, 0.69268, 
    0.68869, 0.68472, 0.68076, 0.67683, 0.67291, 0.669, 0.66512, 0.66126, 
    0.65742, 0.6536, 0.6498, 0.64602, 0.64226, 0.63853, 0.63482, 0.63113, 
    0.62746, 0.62381, 0.62019, 0.6166, 0.61303, 0.60948, 0.60596, 0.60246, 
    0.59899, 0.59554, 0.59212, 0.58873, 0.58536, 0.58201, 0.57869, 0.57539, 
    0.57212, 0.56887, 0.56565, 0.56244, 0.55926, 0.5561, 0.55297, 0.54985, 
    0.54675, 0.54368, 0.54063, 0.53759, 0.53458, 0.53158, 0.52861, 0.52565, 
    0.52272, 0.5198, 0.51691, 0.51403, 0.51117, 0.50833, 0.5055, 0.5027, 
    0.49991, 0.49714, 0.49439, 0.49165, 0.48892, 0.48622, 0.48353, 0.48085, 
    0.47818, 0.47554, 0.4729, 0.47028, 0.46767, 0.46508, 0.4625, 0.45994, 
    0.45739, 0.45485, 0.45233, 0.44982, 0.44733, 0.44485, 0.44239, 0.43994, 
    0.43751, 0.43509, 0.43268, 0.43029, 0.42792, 0.42556, 0.42322, 0.42089, 
    0.41858, 0.41628, 0.414, 0.41174, 0.40949, 0.40726, 0.40504, 0.40284, 
    0.40066, 0.39849, 0.39634, 0.39421, 0.39209, 0.38999, 0.3879, 0.38583, 
    0.38377, 0.38173, 0.3797, 0.37769, 0.37569, 0.3737, 0.37172, 0.36976, 
    0.36781, 0.36587, 0.36394, 0.36203, 0.36012, 0.35823, 0.35635, 0.35448, 
    0.35262, 0.35077, 0.34893, 0.3471, 0.34529, 0.34348, 0.34168, 0.3399, 
    0.33812, 0.33636, 0.33461, 0.33286, 0.33113, 0.32941, 0.3277, 0.326, 
    0.32431, 0.32263, 0.32096, 0.31931, 0.31767, 0.31604, 0.31442, 0.31281, 
    0.31121, 0.30963, 0.30805, 0.30649, 0.30494, 0.3034, 0.30187, 0.30035, 
    0.29883, 0.29733, 0.29583, 0.29434, 0.29285, 0.29138, 0.2899, 0.28844, 
    0.28698, 0.28552, 0.28407, 0.28262, 0.28118, 0.27974, 0.27831, 0.27689, 
    0.27548, 0.27407, 0.27267, 0.27127, 0.26989, 0.26852, 0.26716, 0.26581, 
    0.26447, 0.26315, 0.26183, 0.26053, 0.25925, 0.25797, 0.25671, 0.25546, 
    0.25422, 0.253, 0.25178, 0.25058, 0.24938, 0.2482, 0.24702, 0.24585, 
    0.24469, 0.24354, 0.24239, 0.24125, 0.24012, 0.23899, 0.23787, 0.23675, 
    0.23564, 0.23453, 0.23343, 0.23233, 0.23124, 0.23014, 0.22906, 0.22797, 
    0.22689, 0.22581, 0.22474, 0.22367, 0.22261, 0.22154, 0.22049, 0.21943, 
    0.21839, 0.21734, 0.21631, 0.21527, 0.21425, 0.21323, 0.21221, 0.21121, 
    0.21021, 0.20921, 0.20823, 0.20725, 0.20628, 0.20532, 0.20437, 0.20343, 
    0.20249, 0.20156, 0.20064, 0.19973, 0.19883, 0.19793, 0.19704, 0.19616, 
    0.19529, 0.19442, 0.19356, 0.1927, 0.19186, 0.19101, 0.19018, 0.18935, 
    0.18852, 0.18771, 0.18689, 0.18609, 0.18529, 0.18449, 0.18371, 0.18292, 
    0.18215, 0.18138, 0.18062, 0.17986, 0.17911, 0.17836, 0.17762, 0.17689, 
    0.17616, 0.17544, 0.17473, 0.17402, 0.17332, 0.17263, 0.17195, 0.17128, 
    0.17062, 0.16996, 0.16929, 0.16863, 0.16797, 0.16732, 0.16666, 0.16601, 
    0.16536, 0.16471, 0.16406, 0.16342, 0.16278, 0.16214, 0.1615, 0.16087, 
    0.16024, 0.15961, 0.15898, 0.15836, 0.15774, 0.15712, 0.15651, 0.15589, 
    0.15529, 0.15468, 0.15408, 0.15347, 0.15288, 0.15228, 0.15169, 0.1511, 
    0.15051, 0.14992, 0.14933, 0.14875, 0.14817, 0.14759, 0.14702, 0.14645, 
    0.14588, 0.14531, 0.14474, 0.14418, 0.14362, 0.14306, 0.14251, 0.14195, 
    0.14141, 0.14086, 0.14032, 0.13978, 0.13924, 0.1387, 0.13817, 0.13764, 
    0.13711, 0.13659, 0.13606, 0.13554, 0.13502, 0.1345, 0.13399, 0.13348, 
    0.13296, 0.13245, 0.13194, 0.13144, 0.13093, 0.13043, 0.12993, 0.12943, 
    0.12894, 0.12844, 0.12795, 0.12746, 0.12698, 0.12649, 0.12601, 0.12553, 
    0.12506, 0.12458, 0.12411, 0.12364, 0.12317, 0.12271, 0.12225, 0.12178, 
    0.12132, 0.12087, 0.12041, 0.11995, 0.1195, 0.11905, 0.1186, 0.11815, 
    0.1177, 0.11725, 0.11681, 0.11636, 0.11592, 0.11548, 0.11504, 0.1146, 
    0.11416, 0.11373, 0.11329, 0.11286, 0.11243, 0.112, 0.11157, 0.11114, 
    0.11071, 0.11029, 0.10986, 0.10944, 0.10902, 0.10859, 0.10817, 0.10775, 
    0.10733, 0.10691, 0.1065, 0.10608, 0.10567, 0.10526, 0.10484, 0.10444, 
    0.10403, 0.10362, 0.10322, 0.10282, 0.10242, 0.10202, 0.10162, 0.10123, 
    0.10083, 0.10044, 0.10005, 0.09966, 0.099272, 0.098886, 0.098501, 
    0.098117, 0.097735, 0.097354, 0.096974, 0.096595, 0.096218, 0.095841, 
    0.095466, 0.095092, 0.09472, 0.094348, 0.093978, 0.093609, 0.093242, 
    0.092875, 0.09251, 0.092146, 0.091784, 0.091422, 0.091062, 0.090704, 
    0.090346, 0.08999, 0.089635, 0.089281, 0.088928, 0.088577, 0.088227, 
    0.087878, 0.08753, 0.087184, 0.086839, 0.086495, 0.086153, 0.085812, 
    0.085472, 0.085133, 0.084796, 0.084461, 0.084126, 0.083793, 0.083462, 
    0.083131, 0.082803, 0.082475, 0.082149, 0.081825, 0.081501, 0.081179, 
    0.080858, 0.080539, 0.08022, 0.079903, 0.079586, 0.079271, 0.078956, 
    0.078642, 0.078328, 0.078015, 0.077703, 0.077391, 0.077079, 0.076768, 
    0.076457, 0.076146, 0.075835, 0.075525, 0.075215, 0.074906, 0.074597, 
    0.074289, 0.073981, 0.073674, 0.073368, 0.073064, 0.07276, 0.072457, 
    0.072156, 0.071856, 0.071557, 0.07126, 0.070965, 0.070671, 0.070378, 
    0.070087, 0.069798, 0.069509, 0.069223, 0.068937, 0.068653, 0.06837, 
    0.068088, 0.067807, 0.067527, 0.067248, 0.066969, 0.066692, 0.066416, 
    0.06614, 0.065865, 0.065591, 0.065317, 0.065044, 0.064772, 0.064501, 
    0.06423, 0.06396, 0.06369, 0.063422, 0.063154, 0.062887, 0.06262, 
    0.062354, 0.062089, 0.061825, 0.061561, 0.061298, 0.061036, 0.060774, 
    0.060513, 0.060253, 0.059993, 0.059734, 0.059476, 0.059217, 0.05896, 
    0.058703, 0.058446, 0.05819, 0.057934, 0.057678, 0.057423, 0.057168, 
    0.056913, 0.056658, 0.056404, 0.05615, 0.055896, 0.055642, 0.055388, 
    0.055134, 0.05488, 0.054626, 0.054372, 0.054117, 0.053863, 0.053607, 
    0.053351 ;

 refrac_sigma =
  1.7351, 1.7326, 1.7299, 1.727, 1.7241, 1.721, 1.7181, 1.7152, 1.7124, 
    1.7097, 1.7071, 1.7048, 1.7027, 1.7008, 1.6991, 1.6975, 1.6964, 1.6954, 
    1.6948, 1.6945, 1.6944, 1.6949, 1.6956, 1.697, 1.6988, 1.7011, 1.7041, 
    1.7074, 1.7113, 1.7156, 1.7203, 1.7255, 1.7308, 1.7367, 1.7427, 1.7489, 
    1.7553, 1.7617, 1.7681, 1.7743, 1.7805, 1.7863, 1.7921, 1.7973, 1.8025, 
    1.8074, 1.8121, 1.8166, 1.821, 1.8253, 1.8296, 1.8339, 1.8382, 1.8425, 
    1.8467, 1.851, 1.8553, 1.8595, 1.8637, 1.8679, 1.8721, 1.8762, 1.8802, 
    1.8841, 1.888, 1.8917, 1.8955, 1.8992, 1.903, 1.9068, 1.9106, 1.9144, 
    1.9183, 1.9221, 1.926, 1.9297, 1.9335, 1.9372, 1.9408, 1.9443, 1.9478, 
    1.9512, 1.9545, 1.9577, 1.9609, 1.964, 1.967, 1.97, 1.9728, 1.9755, 
    1.9781, 1.9805, 1.9828, 1.9849, 1.9868, 1.9886, 1.9902, 1.9916, 1.9928, 
    1.9938, 1.9946, 1.9952, 1.9956, 1.9957, 1.9957, 1.9953, 1.9948, 1.9938, 
    1.9926, 1.9911, 1.9893, 1.9873, 1.9851, 1.9827, 1.9802, 1.9778, 1.9753, 
    1.9729, 1.9706, 1.9683, 1.9662, 1.9642, 1.9624, 1.9607, 1.9592, 1.9578, 
    1.9564, 1.9553, 1.9541, 1.9531, 1.9522, 1.9514, 1.9507, 1.9501, 1.9495, 
    1.9491, 1.9487, 1.9484, 1.9481, 1.948, 1.948, 1.948, 1.9481, 1.9482, 
    1.9484, 1.9485, 1.9486, 1.9487, 1.9486, 1.9483, 1.9479, 1.947, 1.9457, 
    1.9441, 1.9414, 1.9383, 1.9343, 1.9293, 1.9237, 1.9165, 1.9087, 1.8995, 
    1.8892, 1.878, 1.8652, 1.8517, 1.8367, 1.8208, 1.804, 1.7859, 1.7673, 
    1.7477, 1.7276, 1.707, 1.686, 1.6647, 1.6434, 1.6222, 1.6012, 1.5807, 
    1.5603, 1.5409, 1.5218, 1.5035, 1.4863, 1.4693, 1.4542, 1.4396, 1.4263, 
    1.4144, 1.4034, 1.3946, 1.3865, 1.38, 1.3748, 1.3704, 1.3676, 1.3653, 
    1.364, 1.3632, 1.3628, 1.3628, 1.3628, 1.3627, 1.3625, 1.3621, 1.3611, 
    1.3599, 1.358, 1.3558, 1.353, 1.3498, 1.3462, 1.3421, 1.3379, 1.3334, 
    1.3286, 1.3238, 1.3187, 1.3136, 1.3084, 1.3032, 1.298, 1.2928, 1.2875, 
    1.2823, 1.2772, 1.2722, 1.2674, 1.2627, 1.2583, 1.2542, 1.2503, 1.2469, 
    1.2437, 1.2409, 1.2384, 1.2361, 1.2343, 1.2326, 1.2313, 1.2301, 1.2291, 
    1.2283, 1.2276, 1.2271, 1.2267, 1.2264, 1.2262, 1.226, 1.2259, 1.2258, 
    1.2257, 1.2257, 1.2257, 1.2257, 1.2257, 1.2258, 1.2258, 1.2258, 1.2258, 
    1.2258, 1.2258, 1.2258, 1.2257, 1.2256, 1.2256, 1.2254, 1.2253, 1.2252, 
    1.2251, 1.225, 1.2248, 1.2247, 1.2246, 1.2245, 1.2244, 1.2243, 1.2243, 
    1.2242, 1.2242, 1.2241, 1.224, 1.224, 1.2239, 1.2239, 1.2239, 1.2238, 
    1.2238, 1.2237, 1.2237, 1.2236, 1.2235, 1.2235, 1.2234, 1.2233, 1.2233, 
    1.2232, 1.2231, 1.223, 1.2229, 1.2228, 1.2227, 1.2225, 1.2224, 1.2222, 
    1.222, 1.2218, 1.2216, 1.2213, 1.2211, 1.2208, 1.2204, 1.2201, 1.2198, 
    1.2194, 1.2191, 1.2187, 1.2183, 1.218, 1.2176, 1.2173, 1.2169, 1.2166, 
    1.2163, 1.2159, 1.2156, 1.2154, 1.2151, 1.2148, 1.2146, 1.2143, 1.2141, 
    1.2139, 1.2137, 1.2135, 1.2134, 1.2132, 1.2131, 1.213, 1.2129, 1.2129, 
    1.2128, 1.2128, 1.2128, 1.2128, 1.2128, 1.2128, 1.2128, 1.2128, 1.2128, 
    1.2128, 1.2127, 1.2127, 1.2126, 1.2124, 1.2123, 1.2121, 1.2119, 1.2116, 
    1.2113, 1.2109, 1.2105, 1.2101, 1.2096, 1.209, 1.2084, 1.2078, 1.2071, 
    1.2063, 1.2055, 1.2047, 1.2038, 1.2029, 1.202, 1.2011, 1.2001, 1.1992, 
    1.1983, 1.1975, 1.1968, 1.1962, 1.1957, 1.1954, 1.1951, 1.195, 1.195, 
    1.195, 1.195, 1.1949, 1.1949, 1.1947, 1.1944, 1.1939, 1.1933, 1.1926, 
    1.1916, 1.1904, 1.1889, 1.1871, 1.185, 1.1824, 1.1796, 1.176, 1.1722, 
    1.1678, 1.1627, 1.1573, 1.1509, 1.1443, 1.137, 1.1292, 1.1211, 1.1122, 
    1.1029, 1.0932, 1.083, 1.0725, 1.0617, 1.0508, 1.0398, 1.0288, 1.0179, 
    1.0074, 0.997, 0.98706, 0.97736, 0.96789, 0.95878, 0.94974, 0.94094, 
    0.93213, 0.92331, 0.9144, 0.9054, 0.89631, 0.88715, 0.87794, 0.86867, 
    0.85932, 0.84997, 0.84056, 0.83112, 0.8217, 0.81224, 0.803, 0.79373, 
    0.7845, 0.77514, 0.76565, 0.75594, 0.74609, 0.73606, 0.72587, 0.71552, 
    0.70516, 0.6947, 0.68422, 0.67366, 0.663, 0.65235, 0.64161, 0.63089, 
    0.62013, 0.60932, 0.5986, 0.58781, 0.5772, 0.56667, 0.55626, 0.54628, 
    0.53638, 0.52711, 0.51806, 0.50937, 0.50121, 0.49322, 0.48602, 0.47907, 
    0.4726, 0.46663, 0.46084, 0.45569, 0.45067, 0.44598, 0.44157, 0.4373, 
    0.4335, 0.42981, 0.42643, 0.42325, 0.4202, 0.41741, 0.41466, 0.41198, 
    0.40932, 0.40667, 0.40397, 0.40124, 0.39843, 0.39554, 0.39257, 0.38947, 
    0.38629, 0.38296, 0.37952, 0.37597, 0.37227, 0.36848, 0.36454, 0.3605, 
    0.35636, 0.35209, 0.34775, 0.34323, 0.33857, 0.33372, 0.32859, 0.32329, 
    0.31754, 0.31156, 0.30517, 0.29842, 0.29139, 0.28394, 0.27626, 0.26828, 
    0.26007, 0.25162, 0.2431, 0.23441, 0.22576, 0.21721, 0.20868, 0.20074, 
    0.19286, 0.18568, 0.17887, 0.17241, 0.16669, 0.16115, 0.15636, 0.15189, 
    0.14781, 0.14428, 0.14092, 0.13809, 0.13545, 0.13309, 0.13103, 0.12909, 
    0.12751, 0.12606, 0.12484, 0.1239, 0.12309, 0.12267, 0.12236, 0.12228, 
    0.12236, 0.12252, 0.12278, 0.12305, 0.12333, 0.12358, 0.12382, 0.124, 
    0.12415, 0.12426, 0.12433, 0.12439, 0.12443, 0.12448, 0.12455, 0.12464, 
    0.12474, 0.12489, 0.12505, 0.12526, 0.12551, 0.1258, 0.12617, 0.12657, 
    0.12705, 0.12756, 0.12812, 0.12872, 0.12933, 0.12994, 0.13054, 0.13111, 
    0.1316, 0.13206, 0.13236, 0.1326, 0.13271, 0.13269, 0.1326, 0.13235, 
    0.13205, 0.13165, 0.1312, 0.13071, 0.13016, 0.1296, 0.12901, 0.12842, 
    0.12782, 0.12723, 0.12663, 0.12602, 0.1254, 0.12478, 0.12416, 0.12354, 
    0.12291, 0.12229, 0.12166, 0.12104, 0.12042, 0.11983, 0.11927, 0.11874, 
    0.11828, 0.11784, 0.11749, 0.11718, 0.11694, 0.11675, 0.1166, 0.11651, 
    0.11643, 0.11637, 0.1163, 0.11623, 0.11613, 0.11602, 0.1159, 0.11576, 
    0.11561, 0.11545, 0.11528, 0.1151, 0.11492, 0.11474, 0.11455, 0.11436, 
    0.11418, 0.11402, 0.11387, 0.11374, 0.11362, 0.11351, 0.11341, 0.11333, 
    0.11326, 0.11319, 0.11314, 0.11308, 0.11303, 0.11299, 0.11295, 0.11292, 
    0.11289, 0.11287, 0.11287, 0.11286, 0.11287, 0.11288, 0.11291, 0.11293, 
    0.11296, 0.11297, 0.11297, 0.11295, 0.1129, 0.11284, 0.11272, 0.11258, 
    0.1124, 0.11219, 0.11196, 0.11171, 0.11145, 0.11118, 0.11091, 0.11063, 
    0.11035, 0.11007, 0.10979, 0.10952, 0.10925, 0.10899, 0.10873, 0.10848, 
    0.10822, 0.10794, 0.10766, 0.10737, 0.10707, 0.10678, 0.10648, 0.1062, 
    0.10592, 0.10565, 0.10539, 0.10515, 0.10493, 0.10474, 0.10459, 0.10446, 
    0.10436, 0.10429, 0.10424, 0.10421, 0.10419, 0.10419, 0.10419, 0.10421, 
    0.10423, 0.10425, 0.10426, 0.10428, 0.10429, 0.10429, 0.10429, 0.10428, 
    0.10426, 0.10425, 0.10423, 0.10422, 0.10421, 0.10421, 0.10421, 0.10424, 
    0.10427, 0.10432, 0.10437, 0.10444, 0.10451, 0.10459, 0.10467, 0.10475, 
    0.10484, 0.10492, 0.105, 0.10509, 0.10517, 0.10524, 0.10531, 0.10538, 
    0.10545, 0.10552, 0.10559, 0.10566, 0.10573, 0.1058, 0.10587, 0.10594, 
    0.106, 0.10607, 0.10613, 0.1062, 0.10626, 0.10632, 0.10638, 0.10643, 
    0.10649, 0.10654, 0.1066, 0.10667, 0.10673, 0.1068, 0.10688, 0.10696, 
    0.10704, 0.10713, 0.10722, 0.10731, 0.10741, 0.10751, 0.10762, 0.10772, 
    0.10783, 0.10794, 0.10806, 0.10817, 0.10828, 0.10839, 0.10849, 0.10859, 
    0.10869, 0.10878, 0.10885, 0.10893, 0.10899, 0.10904, 0.10909, 0.10911, 
    0.10913, 0.10912, 0.10909, 0.10905, 0.10899, 0.10892, 0.10881, 0.10869, 
    0.10854, 0.10835, 0.10814, 0.10789, 0.10762, 0.10733, 0.107, 0.10666, 
    0.10628, 0.10589, 0.10547, 0.10503, 0.10459, 0.10412, 0.10364, 0.10315, 
    0.10264, 0.10213, 0.10159, 0.10106, 0.10052, 0.099987, 0.099449, 
    0.098902, 0.098347, 0.097773, 0.097184, 0.09658, 0.095958, 0.095328, 
    0.094688, 0.094046, 0.093403, 0.092776, 0.092156, 0.091578, 0.091029, 
    0.090521, 0.090075, 0.089654, 0.089308, 0.088989, 0.088717, 0.088488, 
    0.088279, 0.08812, 0.087974, 0.087856, 0.087758, 0.087672, 0.087609, 
    0.087553, 0.087513, 0.087485, 0.087464, 0.087457, 0.087454, 0.087458, 
    0.087465, 0.087475, 0.087489, 0.087504, 0.087523, 0.087542, 0.087562, 
    0.087581, 0.087599, 0.087613, 0.087625, 0.087634, 0.087637, 0.087639, 
    0.087639, 0.087637, 0.087636, 0.087637, 0.087638, 0.087643, 0.087649, 
    0.087659, 0.087669, 0.087679, 0.087689, 0.0877, 0.087709, 0.087719, 
    0.087728, 0.087736, 0.087744, 0.08775, 0.087756, 0.087761, 0.087765, 
    0.087769, 0.087771, 0.087773, 0.087774, 0.087772, 0.087768, 0.08776, 
    0.087748, 0.087732, 0.087708, 0.087682, 0.087647, 0.087609, 0.087567, 
    0.08752, 0.087471, 0.087418, 0.087366, 0.087313, 0.087261, 0.087209, 
    0.087159, 0.08711, 0.087063, 0.087017, 0.086972, 0.086926, 0.08688, 
    0.086831, 0.086777, 0.08672, 0.08665, 0.086574, 0.086482, 0.08637, 
    0.086244, 0.086074, 0.085884, 0.085649, 0.085379, 0.085081, 0.084736, 
    0.084375, 0.083983, 0.083582, 0.083172, 0.082764, 0.082356, 0.08196, 
    0.081576, 0.081204, 0.080855, 0.080514, 0.080189, 0.079865, 0.079544, 
    0.079217, 0.078887, 0.078534, 0.07816, 0.077751, 0.077272, 0.076759, 
    0.076108, 0.075401, 0.074587, 0.07367, 0.072691, 0.071588, 0.070443, 
    0.069222, 0.067972, 0.066693, 0.065464, 0.064256, 0.063149, 0.062149, 
    0.061233, 0.060529, 0.059891, 0.059422, 0.059037, 0.058731, 0.058527, 
    0.058356, 0.058257, 0.058183, 0.058137, 0.058114, 0.058099, 0.058098, 
    0.0581, 0.058107, 0.058119, 0.058132, 0.058152, 0.058178, 0.058212, 
    0.058261, 0.058317, 0.058391, 0.058463, 0.058529, 0.058571, 0.058599, 
    0.058564, 0.058505, 0.058388, 0.058222, 0.058024, 0.057765, 0.057491, 
    0.057188, 0.056884, 0.056579, 0.056309, 0.056057, 0.055858, 0.055689, 
    0.055549, 0.05545, 0.055365, 0.055313, 0.055276, 0.055254, 0.055248, 
    0.055248, 0.055258, 0.05527, 0.055285, 0.055301, 0.055316, 0.05533, 
    0.055344, 0.055358, 0.055372, 0.055386, 0.0554, 0.055412, 0.055421, 
    0.055426, 0.055429, 0.055427, 0.055423, 0.055419, 0.055415, 0.055412, 
    0.055412, 0.055413, 0.055421, 0.055434, 0.055453, 0.055482, 0.055514, 
    0.055556, 0.055603, 0.055656, 0.055718, 0.055783, 0.055858, 0.05594, 
    0.056028, 0.056123, 0.056221, 0.056325, 0.056431, 0.056543, 0.056662, 
    0.056784, 0.056918, 0.057055, 0.057199, 0.057349, 0.057501, 0.057657, 
    0.057815, 0.057976, 0.058141, 0.058307, 0.058477, 0.058647, 0.058818, 
    0.058983, 0.059144, 0.059294, 0.059442, 0.059585, 0.059728, 0.059871, 
    0.060008, 0.060143, 0.060268, 0.060385, 0.060495, 0.060597, 0.060695, 
    0.060792, 0.060888, 0.060982, 0.061067, 0.061149, 0.061224, 0.061298, 
    0.06137, 0.06144, 0.06151, 0.061582, 0.061656, 0.061733, 0.061814, 
    0.061896, 0.06198, 0.062066, 0.062152, 0.062236, 0.062317, 0.062385, 
    0.06245, 0.062506, 0.062557, 0.062604, 0.062645, 0.062684, 0.062718, 
    0.062744, 0.062763, 0.062768, 0.062769, 0.06276, 0.062749, 0.062738, 
    0.062729, 0.06272, 0.06271, 0.062698, 0.062683, 0.062667, 0.062652, 
    0.062645, 0.062644, 0.062648, 0.06266, 0.062676, 0.0627, 0.062724, 
    0.062749, 0.062771, 0.062793, 0.062812, 0.062832, 0.062851, 0.062868, 
    0.062884, 0.062893, 0.062898, 0.062896, 0.06288, 0.062856, 0.062813, 
    0.062767, 0.062714, 0.062653, 0.062586, 0.0625, 0.062409, 0.062304, 
    0.062193, 0.062077, 0.061951, 0.061822, 0.06169, 0.061558, 0.061426, 
    0.061295, 0.061164, 0.061036, 0.060911, 0.060791, 0.060679, 0.060572, 
    0.060477, 0.060389, 0.060313, 0.060253, 0.060201, 0.060163, 0.06013, 
    0.060105, 0.060087, 0.060073, 0.06007, 0.06007, 0.060077, 0.060093, 
    0.060114, 0.060152, 0.060195, 0.060251, 0.060314, 0.060382, 0.060461, 
    0.060543, 0.060634, 0.060727, 0.060822, 0.060916, 0.061008, 0.061096, 
    0.061179, 0.061256, 0.06132, 0.061381, 0.061429, 0.06147, 0.061503, 
    0.061522, 0.061537, 0.06154, 0.06154, 0.061536, 0.061529, 0.061521, 
    0.06151, 0.061499, 0.061487, 0.061477, 0.061467, 0.061461, 0.061456, 
    0.061453, 0.061453, 0.061454, 0.061458, 0.061462, 0.061468, 0.061476, 
    0.061484, 0.061494, 0.061505, 0.061516, 0.061529, 0.061541, 0.061555, 
    0.061568, 0.061582, 0.061596, 0.061611, 0.061627, 0.061642, 0.061657, 
    0.061672, 0.061685, 0.061699, 0.061712, 0.061725, 0.061739, 0.061755, 
    0.061777, 0.061803, 0.061842, 0.061888, 0.061945, 0.062015, 0.062091, 
    0.062183, 0.062277, 0.062379, 0.062484, 0.062591, 0.062705, 0.062821, 
    0.062939, 0.06306, 0.063182, 0.063305, 0.063428, 0.063554, 0.063682, 
    0.063813, 0.06395, 0.06409, 0.064237, 0.064388, 0.064542, 0.064703, 
    0.064865, 0.065037, 0.065214, 0.0654, 0.065595, 0.065793, 0.066, 
    0.066212, 0.066431, 0.066653, 0.066875, 0.067093, 0.067306, 0.06751, 
    0.067702, 0.067888, 0.068056, 0.06822, 0.068376, 0.068527, 0.068675, 
    0.068814, 0.06895, 0.069082, 0.069211, 0.069339, 0.069465, 0.06959, 
    0.069715, 0.069839, 0.069962, 0.070082, 0.070201, 0.070316, 0.07043, 
    0.070544, 0.070659, 0.070775, 0.070891, 0.071007, 0.071121, 0.071235, 
    0.071348, 0.071461, 0.071574, 0.071686, 0.071797, 0.071908, 0.072016, 
    0.072123, 0.072228, 0.072331, 0.072433, 0.072533, 0.072632, 0.07273, 
    0.072825, 0.072919, 0.073007, 0.073094, 0.073176, 0.073254, 0.073329, 
    0.073396, 0.073459, 0.073514, 0.073563, 0.073606, 0.073638, 0.073666, 
    0.073683, 0.073696, 0.073703, 0.073703, 0.073699, 0.073684, 0.073664, 
    0.073635, 0.073598, 0.073557, 0.073506, 0.073452, 0.073394, 0.073331, 
    0.073266, 0.073199, 0.07313, 0.073061, 0.072992, 0.072924, 0.072858, 
    0.072793, 0.072733, 0.072676, 0.072621, 0.072574, 0.072532, 0.072499, 
    0.072475, 0.072457, 0.072449, 0.072446, 0.072452, 0.072465, 0.072482, 
    0.072508, 0.072536, 0.07257, 0.072604, 0.072641, 0.072676, 0.07271, 
    0.072743, 0.072774, 0.072804, 0.072833, 0.072861, 0.072888, 0.072912, 
    0.072935, 0.072953, 0.07297, 0.072981, 0.072989, 0.072994, 0.072996, 
    0.072996, 0.072992, 0.072985, 0.072974, 0.072959, 0.072942, 0.072919, 
    0.072895, 0.072869, 0.072841, 0.072812, 0.07278, 0.072747, 0.072711, 
    0.072674, 0.072635, 0.072593, 0.072551, 0.072507, 0.072462, 0.072415, 
    0.072365, 0.072313, 0.072258, 0.0722, 0.072139, 0.072074, 0.072007, 
    0.071934, 0.071858, 0.071778, 0.071692, 0.071603, 0.071511, 0.071418, 
    0.071323, 0.071226, 0.071127, 0.071025, 0.070923, 0.070819, 0.070716, 
    0.070612, 0.070508, 0.070402, 0.070294, 0.070181, 0.070064, 0.069942, 
    0.069818, 0.069693, 0.069565, 0.069434, 0.069299, 0.069162, 0.069019, 
    0.068871, 0.068717, 0.068557, 0.068393, 0.068221, 0.068045, 0.067863, 
    0.067677, 0.06749, 0.067303, 0.067114, 0.066926, 0.066738, 0.066551, 
    0.066369, 0.066189, 0.066012, 0.065837, 0.065663, 0.065495, 0.065326, 
    0.065159, 0.06499, 0.064819, 0.064645, 0.06447, 0.064294, 0.064119, 
    0.063943, 0.06377, 0.063598, 0.063429, 0.063263, 0.063099, 0.06294, 
    0.062784, 0.062639, 0.0625, 0.06237, 0.062253, 0.06214, 0.062042, 
    0.061951, 0.061869, 0.0618, 0.061736, 0.061683, 0.061632, 0.061586, 
    0.061544, 0.061502, 0.061462, 0.061419, 0.061372, 0.061319, 0.061264, 
    0.061198, 0.061126, 0.061044, 0.060955, 0.060862, 0.060762, 0.060661, 
    0.060554, 0.060444, 0.06033, 0.060212, 0.060092, 0.05997, 0.059848, 
    0.059725, 0.059607, 0.059491, 0.059379, 0.059267, 0.059156, 0.059048, 
    0.058941, 0.05884, 0.058742, 0.058648, 0.058559, 0.058473, 0.0584, 
    0.058332, 0.058272, 0.058221, 0.058173, 0.058142, 0.058118, 0.058107, 
    0.058109, 0.058116, 0.058141, 0.058172, 0.058218, 0.058276, 0.05834, 
    0.058419, 0.058504, 0.058603, 0.058716, 0.058839, 0.058985, 0.05914, 
    0.059315, 0.0595, 0.059695, 0.059905, 0.060119, 0.060342, 0.060568, 
    0.060796, 0.061021, 0.061242, 0.061446, 0.06164, 0.061821, 0.061991, 
    0.062155, 0.062301, 0.062437, 0.062555, 0.062657, 0.062751, 0.062827, 
    0.062898, 0.062958, 0.063012, 0.063062, 0.063107, 0.06315, 0.063189, 
    0.063226, 0.063261, 0.063294, 0.063327, 0.063358, 0.063388, 0.063417, 
    0.063444, 0.06347, 0.063493, 0.063513, 0.063532, 0.063547, 0.063561, 
    0.063572, 0.063582, 0.06359, 0.063595, 0.063598, 0.063597, 0.063593, 
    0.063586, 0.063576, 0.063564, 0.063547, 0.063528, 0.063506, 0.06348, 
    0.063453, 0.063422, 0.06339, 0.063356, 0.063322, 0.063288, 0.063251, 
    0.063214, 0.063175, 0.063134, 0.063091, 0.063041, 0.062987, 0.062925, 
    0.062855, 0.062778, 0.062689, 0.062597, 0.062498, 0.062399, 0.062298, 
    0.062197, 0.062095, 0.061994, 0.061892, 0.061789, 0.061685, 0.061579, 
    0.061469, 0.061356, 0.061239, 0.061112, 0.060982, 0.060839, 0.060691, 
    0.060534, 0.060371, 0.060203, 0.060028, 0.059849, 0.059664, 0.059469, 
    0.05927, 0.059063, 0.058853, 0.058639, 0.058418, 0.058193, 0.057969, 
    0.057747, 0.057532, 0.057327, 0.057131, 0.056955, 0.056786, 0.056634, 
    0.056487, 0.056346, 0.056209, 0.056074, 0.05594, 0.055806, 0.05567, 
    0.055531, 0.055389, 0.055241, 0.05509, 0.054936, 0.054779, 0.054622, 
    0.054466, 0.054312, 0.05416, 0.05401, 0.053861, 0.053711, 0.053562, 
    0.053414, 0.053269, 0.053126, 0.052989, 0.052854, 0.052723, 0.052597, 
    0.052472, 0.052358, 0.052246, 0.052142, 0.052044, 0.051952, 0.051866, 
    0.051783, 0.051705, 0.051627, 0.051549, 0.051471, 0.051393, 0.051314, 
    0.051233, 0.051152, 0.051069, 0.050987, 0.050904, 0.050823, 0.050744, 
    0.050668, 0.050594, 0.050526, 0.050461, 0.050399, 0.050341, 0.050285, 
    0.050233, 0.050185, 0.05014, 0.050099, 0.05006, 0.050026, 0.049993, 
    0.049963, 0.049935, 0.049907, 0.049881, 0.049857, 0.049833, 0.049811, 
    0.049791, 0.049772, 0.049754, 0.049736, 0.049719, 0.049701, 0.049684, 
    0.049667, 0.04965, 0.049633, 0.049615, 0.049596, 0.049577, 0.049557, 
    0.049536, 0.049516, 0.049494, 0.049473, 0.049452, 0.049432, 0.049412, 
    0.049395, 0.049379, 0.049369, 0.049362, 0.049361, 0.049364, 0.049369, 
    0.049378, 0.049389, 0.049402, 0.049418, 0.049434, 0.049456, 0.049479, 
    0.049503, 0.049526, 0.049548, 0.049563, 0.049576, 0.049584, 0.049592, 
    0.049599, 0.049605, 0.049611, 0.049615, 0.049617, 0.049619, 0.049619, 
    0.049619, 0.04962, 0.049621, 0.049623, 0.049626, 0.049629, 0.049633, 
    0.049636, 0.049638, 0.049641, 0.049643, 0.049645, 0.049646, 0.049648, 
    0.049647, 0.049646, 0.049642, 0.049638, 0.049633, 0.049628, 0.049623, 
    0.049618, 0.049611, 0.049602, 0.04959, 0.049576, 0.049561, 0.049549, 
    0.049542, 0.049538, 0.049536, 0.049537, 0.049538, 0.049543, 0.049555, 
    0.049572, 0.049603, 0.049638, 0.049683, 0.049728, 0.049772, 0.049814, 
    0.049854, 0.049893, 0.049934, 0.049975, 0.050018, 0.050061, 0.050104, 
    0.050147, 0.05019, 0.050233, 0.050275, 0.050321, 0.050369, 0.050419, 
    0.050469, 0.050518, 0.050561, 0.050602, 0.050635, 0.050663, 0.050688, 
    0.050708, 0.050726, 0.050742, 0.050756, 0.050769, 0.05078, 0.05079, 
    0.0508, 0.050811, 0.050823, 0.050839, 0.050857, 0.050881, 0.050909, 
    0.050942, 0.050981, 0.051023, 0.051075, 0.051132, 0.051196, 0.051271, 
    0.05135, 0.051448, 0.05155, 0.051661, 0.051776, 0.051894, 0.05201, 
    0.052122, 0.052229, 0.05234, 0.052452, 0.052574, 0.052697, 0.052827, 
    0.052959, 0.053093, 0.053233, 0.053374, 0.053519, 0.053662, 0.053806, 
    0.053948, 0.054087, 0.054219, 0.054343, 0.054457, 0.054555, 0.054645, 
    0.054713, 0.054773, 0.054822, 0.054861, 0.054897, 0.054924, 0.054949, 
    0.054968, 0.054981, 0.054991, 0.054989, 0.054983, 0.05497, 0.054954, 
    0.054936, 0.054911, 0.054883, 0.054849, 0.054807, 0.05476, 0.054696, 
    0.054627, 0.054543, 0.054449, 0.054348, 0.054231, 0.05411, 0.053977, 
    0.053837, 0.053689, 0.053529, 0.053363, 0.05318, 0.052988, 0.052785, 
    0.052563, 0.052332, 0.052076, 0.051808, 0.051524, 0.051221, 0.050908, 
    0.05057, 0.050223, 0.049861, 0.049487, 0.049107, 0.048725, 0.048346, 
    0.047978, 0.04762, 0.047267, 0.046927, 0.046593, 0.046275, 0.045979, 
    0.045696, 0.045452, 0.045218, 0.045013, 0.044826, 0.044653, 0.044506, 
    0.044368, 0.044249, 0.044142, 0.044046, 0.043964, 0.043887, 0.043822, 
    0.043761, 0.043707, 0.043659, 0.043615, 0.043576, 0.04354, 0.043508, 
    0.04348, 0.043454, 0.043431, 0.043409, 0.043389, 0.043371, 0.043354, 
    0.04334, 0.043326, 0.043316, 0.043307, 0.0433, 0.043295, 0.043291, 
    0.043289, 0.043289, 0.043289, 0.043291, 0.043293, 0.043295, 0.043296, 
    0.043296, 0.043295, 0.043293, 0.04329, 0.043286, 0.04328, 0.043272, 
    0.043263, 0.043252, 0.043238, 0.043222, 0.043202, 0.043181, 0.043154, 
    0.043122, 0.043085, 0.043042, 0.042996, 0.042945, 0.042893, 0.042841, 
    0.042792, 0.042744, 0.042707, 0.042674, 0.04265, 0.042635, 0.042625, 
    0.04263, 0.04264, 0.042661, 0.042688, 0.042721, 0.04276, 0.042799, 
    0.04284, 0.042879, 0.042915, 0.042945, 0.042973, 0.042994, 0.04301, 
    0.043021, 0.043023, 0.043022, 0.04301, 0.042994, 0.042972, 0.042942, 
    0.04291, 0.04287, 0.042827, 0.042782, 0.042735, 0.042689, 0.042647, 
    0.042608, 0.042572, 0.042542, 0.042515, 0.042495, 0.042479, 0.042468, 
    0.042461, 0.042457, 0.042458, 0.042459, 0.04246, 0.042461, 0.04246, 
    0.042455, 0.042448, 0.042437, 0.042422, 0.042404, 0.04238, 0.042354, 
    0.042322, 0.042286, 0.042248, 0.042204, 0.042158, 0.042107, 0.042053, 
    0.041995, 0.041932, 0.041867, 0.041797, 0.041726, 0.041653, 0.041583, 
    0.041514, 0.041452, 0.041395, 0.041343, 0.041299, 0.041258, 0.041228, 
    0.041202, 0.041182, 0.041169, 0.041159, 0.041159, 0.041162, 0.041174, 
    0.041193, 0.041216, 0.041248, 0.041284, 0.041326, 0.041372, 0.04142, 
    0.041471, 0.041521, 0.041567, 0.041609, 0.041646, 0.041675, 0.041701, 
    0.04172, 0.041737, 0.041751, 0.041761, 0.041771, 0.041777, 0.041782, 
    0.041786, 0.041788, 0.041789, 0.041787, 0.041783, 0.041777, 0.041767, 
    0.041756, 0.04174, 0.041722, 0.041699, 0.041671, 0.041641, 0.041604, 
    0.041564, 0.041519, 0.041471, 0.04142, 0.041366, 0.041312, 0.041257, 
    0.041201, 0.041143, 0.041085, 0.041027, 0.040968, 0.040909, 0.040851, 
    0.040795, 0.040739, 0.040685, 0.040635, 0.040588, 0.040552, 0.040519, 
    0.0405, 0.040487, 0.040481, 0.040484, 0.040489, 0.040503, 0.040518, 
    0.040538, 0.040561, 0.040586, 0.040613, 0.040639, 0.040665, 0.040692, 
    0.04072, 0.04075, 0.040781, 0.040815, 0.040852, 0.040892, 0.040936, 
    0.040982, 0.041032, 0.041084, 0.041137, 0.041194, 0.041251, 0.041308, 
    0.041365, 0.041422, 0.041478, 0.041534, 0.041591, 0.041649, 0.041707, 
    0.041763, 0.041819, 0.041868, 0.041915, 0.041958, 0.041996, 0.042033, 
    0.042068, 0.042102, 0.042135, 0.042165, 0.042195, 0.042223, 0.042254, 
    0.042289, 0.042333, 0.042381, 0.04244, 0.042502, 0.04257, 0.042641, 
    0.042712, 0.042783, 0.042855, 0.042929, 0.043007, 0.043089, 0.04318, 
    0.043273, 0.043372, 0.043476, 0.043585, 0.043705, 0.043832, 0.043975, 
    0.044127, 0.044289, 0.044463, 0.044639, 0.044823, 0.045008, 0.045194, 
    0.045377, 0.045558, 0.045726, 0.045888, 0.04604, 0.04618, 0.046316, 
    0.046432, 0.046541, 0.046634, 0.046712, 0.046781, 0.046831, 0.046874, 
    0.046902, 0.046915, 0.046918, 0.046892, 0.046854, 0.046787, 0.046701, 
    0.0466, 0.046474, 0.046342, 0.046195, 0.046042, 0.045882, 0.0457, 
    0.04551, 0.045296, 0.045072, 0.044835, 0.044583, 0.044324, 0.044048, 
    0.043764, 0.043471, 0.043173, 0.042873, 0.042576, 0.042283, 0.041998, 
    0.04173, 0.041469, 0.04124, 0.041021, 0.040825, 0.040647, 0.040478, 
    0.040333, 0.040195, 0.040073, 0.039964, 0.039863, 0.039784, 0.039711, 
    0.039655, 0.039609, 0.039572, 0.039546, 0.039525, 0.039513, 0.039504, 
    0.0395, 0.039504, 0.039511, 0.039527, 0.039546, 0.039569, 0.039593, 
    0.039618, 0.039643, 0.039667, 0.039689, 0.03971, 0.039731, 0.039749, 
    0.039766, 0.039781, 0.039792, 0.039801, 0.039805, 0.039808, 0.03981, 
    0.039812, 0.039814, 0.039816, 0.039818, 0.03982, 0.039821, 0.039822, 
    0.039824, 0.039825, 0.039826, 0.039828, 0.039829, 0.03983, 0.039832, 
    0.039833, 0.039835, 0.039838, 0.039841, 0.039844, 0.039848, 0.039852, 
    0.039856, 0.039861, 0.039867, 0.039875, 0.039885, 0.039896, 0.03991, 
    0.039926, 0.039945, 0.039967, 0.039992, 0.040019, 0.040047, 0.040076, 
    0.040105, 0.040133, 0.04016, 0.040187, 0.040213, 0.040237, 0.040259, 
    0.040279, 0.040296, 0.040309, 0.04032, 0.040329, 0.040338, 0.040345, 
    0.040352, 0.040359, 0.040365, 0.040372, 0.040379, 0.040387, 0.040395, 
    0.040405, 0.040417, 0.04043, 0.040446, 0.040462, 0.040478, 0.040495, 
    0.040511, 0.040527, 0.040543, 0.040559, 0.040576, 0.040593, 0.040612, 
    0.040631, 0.040652, 0.040674, 0.040697, 0.040721, 0.040746, 0.040773, 
    0.0408, 0.040828, 0.040856, 0.040884, 0.040911, 0.040938, 0.040962, 
    0.040986, 0.041009, 0.041032, 0.041054, 0.041073, 0.041088, 0.0411, 
    0.041103, 0.041103, 0.041095, 0.041083, 0.041068, 0.041051, 0.041033, 
    0.041015, 0.040995, 0.040975, 0.040955, 0.040934, 0.040915, 0.040895, 
    0.040876, 0.040855, 0.040834, 0.040811, 0.04079, 0.040769, 0.04075, 
    0.040733, 0.040717, 0.040703, 0.040689, 0.040678, 0.040668, 0.040662, 
    0.040658, 0.040657, 0.040658, 0.04066, 0.040664, 0.040669, 0.040675, 
    0.040683, 0.040693, 0.040704, 0.040716, 0.040728, 0.04074, 0.040751, 
    0.040762, 0.040773, 0.040784, 0.040796, 0.040808, 0.040819, 0.04083, 
    0.04084, 0.040851, 0.040863, 0.040877, 0.040893, 0.040912, 0.040933, 
    0.040957, 0.040982, 0.041008, 0.041039, 0.041071, 0.041109, 0.041151, 
    0.041196, 0.041249, 0.041303, 0.041363, 0.041426, 0.041493, 0.041565, 
    0.041637, 0.041708, 0.041775, 0.041838, 0.041891, 0.041941, 0.041984, 
    0.042023, 0.042058, 0.042089, 0.042119, 0.042146, 0.042174, 0.042203, 
    0.042238, 0.042275, 0.04232, 0.042369, 0.042421, 0.042473, 0.042525, 
    0.042575, 0.042624, 0.042671, 0.042717, 0.04276, 0.0428, 0.042838, 
    0.042872, 0.042902, 0.042929, 0.042952, 0.042974, 0.042992, 0.043009, 
    0.043025, 0.04304, 0.043054, 0.043069, 0.043085, 0.043102, 0.04312, 
    0.043139, 0.043158, 0.043177, 0.043196, 0.043215, 0.043234, 0.043253, 
    0.043274, 0.043295, 0.043316, 0.043338, 0.043359, 0.043381, 0.043402, 
    0.043422, 0.043442, 0.043461, 0.043478, 0.043494, 0.043508, 0.043522, 
    0.043532, 0.043543, 0.043554, 0.043565, 0.043577, 0.043592, 0.043608, 
    0.043629, 0.043654, 0.043682, 0.043714, 0.043747, 0.043781, 0.043815, 
    0.043849, 0.043882, 0.043914, 0.043947, 0.043979, 0.04401, 0.044042, 
    0.044073, 0.044104, 0.044134, 0.044166, 0.044196, 0.044227, 0.044256, 
    0.044284, 0.044311, 0.044337, 0.044363, 0.044389, 0.044416, 0.044443, 
    0.044469, 0.044494, 0.044518, 0.044542, 0.044566, 0.044588, 0.04461, 
    0.044623, 0.044634, 0.044635, 0.044628, 0.044615, 0.04459, 0.044562, 
    0.044531, 0.0445, 0.044468, 0.044437, 0.044408, 0.044382, 0.044357, 
    0.044333, 0.04431, 0.044287, 0.044264, 0.044241, 0.044217, 0.04419, 
    0.044162, 0.044127, 0.04409, 0.044048, 0.044002, 0.043953, 0.0439, 
    0.043847, 0.043793, 0.043739, 0.043685, 0.043633, 0.043583, 0.043537, 
    0.043493, 0.043451, 0.043408, 0.043366, 0.043324, 0.043285, 0.043247, 
    0.04321, 0.043173, 0.043133, 0.043092, 0.043049, 0.043003, 0.042958, 
    0.042916, 0.042878, 0.042845, 0.042821, 0.042801, 0.04279, 0.042784, 
    0.042782, 0.042787, 0.042794, 0.04281, 0.042828, 0.04285, 0.042874, 
    0.042899, 0.042923, 0.042947, 0.04297, 0.042992, 0.043014, 0.043033, 
    0.043052, 0.043069, 0.043085, 0.043101, 0.043114, 0.043127, 0.043138, 
    0.04315, 0.043162, 0.043176, 0.04319, 0.043205, 0.043219, 0.043233, 
    0.043243, 0.043252, 0.043258, 0.043262, 0.043265, 0.043265, 0.043264, 
    0.043259, 0.043251, 0.04324, 0.043225, 0.043209, 0.043191, 0.043171, 
    0.043151, 0.043131, 0.043111, 0.043091, 0.04307, 0.04305, 0.043031, 
    0.043013, 0.042997, 0.042981, 0.042966, 0.042954, 0.042942, 0.042936, 
    0.042931, 0.04293, 0.042929, 0.042929, 0.042929, 0.042929, 0.04293, 
    0.042931, 0.042932, 0.042935, 0.042937, 0.042941, 0.042945, 0.042949, 
    0.042954, 0.042959, 0.042965, 0.042972, 0.042978, 0.042985, 0.042992, 
    0.043, 0.043008, 0.043017, 0.043029, 0.043041, 0.043056, 0.043073, 
    0.043092, 0.043112, 0.043132, 0.043152, 0.04317, 0.043186, 0.043198, 
    0.043207, 0.043208, 0.043207, 0.043202, 0.043194, 0.043185, 0.043175, 
    0.043164, 0.043153, 0.043144, 0.043136, 0.043132, 0.04313, 0.043132, 
    0.043135, 0.043139, 0.043145, 0.043152, 0.04316, 0.04317, 0.04318, 
    0.043192, 0.043205, 0.043221, 0.043237, 0.043253, 0.04327, 0.043287, 
    0.043304, 0.043322, 0.043341, 0.043361, 0.043383, 0.043408, 0.043434, 
    0.043462, 0.043492, 0.043523, 0.043559, 0.043596, 0.043638, 0.043683, 
    0.04373, 0.043779, 0.043827, 0.043872, 0.043914, 0.043952, 0.043984, 
    0.044014, 0.044037, 0.044057, 0.044073, 0.044084, 0.044094, 0.0441, 
    0.044106, 0.044111, 0.044117, 0.044124, 0.044134, 0.044144, 0.044156, 
    0.044169, 0.044181, 0.044193, 0.044203, 0.044212, 0.044217, 0.044222, 
    0.044222, 0.044221, 0.044219, 0.044216, 0.044213, 0.044212, 0.044211, 
    0.044212, 0.044214, 0.044216, 0.044219, 0.044222, 0.044225, 0.044227, 
    0.04423, 0.044233, 0.044237, 0.04424, 0.044244, 0.044247, 0.04425, 
    0.044252, 0.044252, 0.044251, 0.044249, 0.044245, 0.044239, 0.044232, 
    0.044225, 0.044218, 0.044211, 0.044204, 0.044197, 0.044189, 0.044181, 
    0.044171, 0.044162, 0.04415, 0.044139, 0.044126, 0.044111, 0.044095, 
    0.044075, 0.044055, 0.044032, 0.044008, 0.043983, 0.043957, 0.043931, 
    0.043902, 0.04387, 0.043836, 0.043797, 0.043755, 0.043709, 0.04366, 
    0.043608, 0.04355, 0.043489, 0.043422, 0.043352, 0.04328, 0.043208, 
    0.043135, 0.043065, 0.042995, 0.042925, 0.042854, 0.042782, 0.04271, 
    0.042638, 0.042566, 0.042496, 0.042426, 0.042359, 0.042291, 0.042224, 
    0.042157, 0.042091, 0.042029, 0.041968, 0.041909, 0.041851, 0.041795, 
    0.04174, 0.041685, 0.041631, 0.04158, 0.04153, 0.041484, 0.04144, 
    0.041399, 0.041361, 0.041324, 0.041291, 0.04126, 0.041232, 0.041206, 
    0.041182, 0.04116, 0.041138, 0.041118, 0.041099, 0.04108, 0.041063, 
    0.041046, 0.041029, 0.041013, 0.040996, 0.040979, 0.04096, 0.040941, 
    0.040922, 0.040901, 0.04088, 0.040858, 0.040834, 0.040809, 0.040783, 
    0.040755, 0.040727, 0.040698, 0.040669, 0.040639, 0.040609, 0.040579, 
    0.040547, 0.040514, 0.04048, 0.040445, 0.040408, 0.040369, 0.040329, 
    0.040287, 0.040245, 0.040202, 0.040159, 0.040116, 0.040072, 0.040026, 
    0.039978, 0.039927, 0.039875, 0.03982, 0.039765, 0.039712, 0.039664, 
    0.039618, 0.039588, 0.039565, 0.039556, 0.039562, 0.039577, 0.039615, 
    0.039661, 0.039725, 0.0398, 0.039884, 0.039974, 0.040064, 0.04015, 
    0.040229, 0.040302, 0.040364, 0.040422, 0.040469, 0.040513, 0.040551, 
    0.040581, 0.040608, 0.040624, 0.040635, 0.040637, 0.040628, 0.040614, 
    0.04059, 0.040562, 0.040529, 0.040492, 0.040453, 0.040404, 0.040351, 
    0.040288, 0.040215, 0.040136, 0.040038, 0.039933, 0.039812, 0.039679, 
    0.039539, 0.039384, 0.039226, 0.039058, 0.038884, 0.038705, 0.038521, 
    0.038337, 0.038153, 0.037975, 0.0378, 0.037636, 0.037476, 0.037326, 
    0.037182, 0.037044, 0.036916, 0.036791, 0.036678, 0.036568, 0.036464, 
    0.036367, 0.036272, 0.036185, 0.036098, 0.036015, 0.035932, 0.035849, 
    0.035765, 0.035681, 0.035596, 0.035511, 0.035426, 0.035343, 0.035261, 
    0.035181, 0.035105, 0.03503, 0.034966, 0.034906, 0.034855, 0.034812, 
    0.034775, 0.034747, 0.034722, 0.034704, 0.034689, 0.034676, 0.034667, 
    0.034659, 0.034653, 0.034648, 0.034644, 0.03464, 0.034635, 0.03463, 
    0.034624, 0.034619, 0.034615, 0.034611, 0.034609, 0.034608, 0.034608, 
    0.034611, 0.034615, 0.034623, 0.034634, 0.034649, 0.034667, 0.034687, 
    0.034712, 0.034738, 0.034767, 0.034799, 0.034832, 0.03487, 0.03491, 
    0.034952, 0.034996, 0.035041, 0.035088, 0.035135, 0.035183, 0.03523, 
    0.035278, 0.035325, 0.035372, 0.035419, 0.035464, 0.035509, 0.035553, 
    0.035597, 0.035641, 0.035685, 0.035728, 0.035768, 0.035808, 0.035845, 
    0.035879, 0.035912, 0.035941, 0.03597, 0.035994, 0.036018, 0.036038, 
    0.036054, 0.036069, 0.036078, 0.036086, 0.036091, 0.036093, 0.036093, 
    0.036087, 0.036079, 0.036066, 0.036047, 0.036026, 0.035999, 0.035971, 
    0.03594, 0.035909, 0.035878, 0.035849, 0.035821, 0.035797, 0.035776, 
    0.035759, 0.035745, 0.035733, 0.035723, 0.035714, 0.035706, 0.035698, 
    0.035689, 0.035681, 0.035672, 0.035663, 0.035654, 0.035645, 0.035636, 
    0.035628, 0.03562, 0.035612, 0.035606, 0.035601, 0.035596, 0.035593, 
    0.035592, 0.035591, 0.035594, 0.035598, 0.035604, 0.035613, 0.035622, 
    0.035633, 0.035644, 0.035654, 0.035664, 0.035673, 0.03568, 0.035687, 
    0.035689, 0.035687, 0.03568, 0.035666, 0.03565, 0.03563, 0.035611, 
    0.035593, 0.035578, 0.035565, 0.035555, 0.035545, 0.035536, 0.035524, 
    0.035511, 0.035496, 0.035479, 0.035461, 0.035441, 0.035421, 0.035401, 
    0.03538, 0.035359, 0.03534, 0.035322, 0.035306, 0.035292, 0.035282, 
    0.035274, 0.035268, 0.035268, 0.03527, 0.035277, 0.035287, 0.0353, 
    0.035319, 0.035339, 0.035365, 0.035394, 0.035427, 0.035466, 0.035508, 
    0.035556, 0.035607, 0.035661, 0.035718, 0.035775, 0.035833, 0.035891, 
    0.035949, 0.036004, 0.036058, 0.036109, 0.036159, 0.036207, 0.036253, 
    0.036299, 0.036345, 0.036391, 0.036438, 0.036485, 0.036531, 0.036576, 
    0.036621, 0.036664, 0.036706, 0.036747, 0.036783, 0.036817, 0.036847, 
    0.036872, 0.036895, 0.036911, 0.036924, 0.036932, 0.036938, 0.036941, 
    0.036943, 0.036946, 0.036948, 0.036951, 0.036955, 0.03696, 0.036966, 
    0.036972, 0.03698, 0.036987, 0.036996, 0.037005, 0.037016, 0.03703, 
    0.037046, 0.037069, 0.037094, 0.037132, 0.037176, 0.037233, 0.037303, 
    0.037382, 0.037483, 0.037592, 0.037717, 0.037853, 0.037998, 0.038156, 
    0.038318, 0.038487, 0.038659, 0.038832, 0.039004, 0.039174, 0.039337, 
    0.039495, 0.039647, 0.03979, 0.03993, 0.040063, 0.040193, 0.040321, 
    0.040446, 0.04057, 0.040692, 0.040813, 0.040934, 0.041055, 0.041175, 
    0.041293, 0.041408, 0.041519, 0.041624, 0.041725, 0.041812, 0.041894, 
    0.041966, 0.042028, 0.042085, 0.04213, 0.042172, 0.042207, 0.042237, 
    0.042264, 0.042286, 0.042307, 0.042326, 0.042342, 0.042357, 0.04237, 
    0.042382, 0.042392, 0.042402, 0.042411, 0.042419, 0.042427, 0.042435, 
    0.042441, 0.042447, 0.042451, 0.042454, 0.042453, 0.042451, 0.042446, 
    0.042439, 0.042431, 0.04242, 0.042408, 0.042396, 0.042382, 0.042368, 
    0.042353, 0.042337, 0.042322, 0.042307, 0.042292, 0.042277, 0.042261, 
    0.042245, 0.042227, 0.042208, 0.042181, 0.042151, 0.04211, 0.042059, 
    0.041999, 0.04192, 0.041833, 0.041725, 0.041607, 0.041475, 0.041329, 
    0.041178, 0.041019, 0.040859, 0.040697, 0.040537, 0.040377, 0.040221, 
    0.040069, 0.039921, 0.039779, 0.039638, 0.039505, 0.039374, 0.039248, 
    0.039126, 0.039007, 0.038893, 0.03878, 0.038669, 0.038556, 0.038441, 
    0.038325, 0.038208, 0.038092, 0.037981, 0.037874, 0.037778, 0.037686, 
    0.037606, 0.037537, 0.037477, 0.037433, 0.037394, 0.037369, 0.037349, 
    0.037334, 0.037324, 0.037315, 0.03731, 0.037305, 0.037302, 0.037299, 
    0.037298, 0.037297, 0.037298, 0.037301, 0.037305, 0.037312, 0.037322, 
    0.037335, 0.037351, 0.037371, 0.037393, 0.037421, 0.03745, 0.037483, 
    0.037518, 0.037556, 0.037596, 0.037637, 0.037679, 0.037721, 0.037765, 
    0.037809, 0.037854, 0.037901, 0.03795, 0.038, 0.038051, 0.038102, 
    0.038152, 0.0382, 0.038247, 0.03829, 0.038332, 0.038368, 0.038401, 
    0.038431, 0.038455, 0.038477, 0.038492, 0.038506, 0.038516, 0.038523, 
    0.038529, 0.038532, 0.038535, 0.038536, 0.038536, 0.038536, 0.038536, 
    0.038535, 0.038534, 0.038534, 0.038534, 0.038534, 0.038534, 0.038534, 
    0.038533, 0.038531, 0.038526, 0.03852, 0.038512, 0.038501, 0.038489, 
    0.038472, 0.038453, 0.038428, 0.038401, 0.038372, 0.038341, 0.038309, 
    0.038277, 0.038246, 0.038215, 0.038184, 0.038155, 0.038127, 0.0381, 
    0.038075, 0.038052, 0.03803, 0.03801, 0.03799, 0.037971, 0.037953, 
    0.037935, 0.037921, 0.037909, 0.037899, 0.037891, 0.037885, 0.037881, 
    0.037879, 0.03788, 0.037883, 0.037887, 0.037895, 0.037905, 0.037917, 
    0.037931, 0.037946, 0.037964, 0.037983, 0.038004, 0.038026, 0.038051, 
    0.038078, 0.038105, 0.038134, 0.038163, 0.038192, 0.03822, 0.038248, 
    0.038275, 0.038301, 0.038326, 0.038349, 0.038372, 0.038393, 0.038414, 
    0.038434, 0.038454, 0.038474, 0.038495, 0.038516, 0.038537, 0.038559, 
    0.038582, 0.038605, 0.038628, 0.038651, 0.038673, 0.038694, 0.038714, 
    0.038733, 0.038751, 0.038766, 0.03878, 0.03879, 0.038798, 0.038802, 
    0.038804, 0.038804, 0.038802, 0.038801, 0.038799, 0.038798, 0.038799, 
    0.038803, 0.038807, 0.038815, 0.038824, 0.038835, 0.038851, 0.038868, 
    0.038891, 0.038916, 0.038945, 0.038976, 0.039008, 0.039041, 0.039075, 
    0.039109, 0.039146, 0.039182, 0.039222, 0.039263, 0.039305, 0.039348, 
    0.039391, 0.03943, 0.039469, 0.039502, 0.039533, 0.03956, 0.039584, 
    0.039605, 0.039623, 0.039638, 0.039651, 0.039661, 0.039671, 0.039678, 
    0.039683, 0.039688, 0.039691, 0.039693, 0.039692, 0.03969, 0.039686, 
    0.039678, 0.039669, 0.039653, 0.039635, 0.039613, 0.039587, 0.039559, 
    0.039528, 0.039497, 0.039464, 0.039432, 0.039399, 0.039368, 0.039339, 
    0.039311, 0.039286, 0.039262, 0.03924, 0.039219, 0.039198, 0.039177, 
    0.039156, 0.039135, 0.039115, 0.039095, 0.039076, 0.039058, 0.039043, 
    0.039028, 0.039017, 0.039009, 0.039004, 0.039004, 0.039007, 0.039016, 
    0.039028, 0.039044, 0.039063, 0.039083, 0.039105, 0.039126, 0.039147, 
    0.039167, 0.039187, 0.039205, 0.039223, 0.039239, 0.039254, 0.039268, 
    0.039281, 0.039292, 0.039302, 0.039309, 0.039315, 0.039313, 0.039309, 
    0.039296, 0.039273, 0.039242, 0.039194, 0.039138, 0.039064, 0.038979, 
    0.038882, 0.038768, 0.038649, 0.038515, 0.038376, 0.03823, 0.038079, 
    0.037927, 0.037774, 0.037623, 0.037475, 0.037335, 0.037199, 0.037073, 
    0.036949, 0.036831, 0.036715, 0.036601, 0.036489, 0.036378, 0.036267, 
    0.036157, 0.036046, 0.035934, 0.035823, 0.035713, 0.035607, 0.035504, 
    0.035411, 0.035322, 0.035246, 0.03518, 0.035122, 0.035079, 0.035042, 
    0.035016, 0.034996, 0.034982, 0.034976, 0.034971, 0.034973, 0.034976, 
    0.034981, 0.034989, 0.034999, 0.035011, 0.035025, 0.03504, 0.035057, 
    0.035074, 0.035093, 0.035112, 0.035132, 0.035152, 0.035173, 0.035196, 
    0.035219, 0.035243, 0.035267, 0.035291, 0.035316, 0.03534, 0.035363, 
    0.035384, 0.035403, 0.03542, 0.035435, 0.035447, 0.035458, 0.035467, 
    0.035474, 0.03548, 0.035484, 0.035487, 0.035488, 0.035487, 0.035485, 
    0.03548, 0.035472, 0.035461, 0.035444, 0.035425, 0.0354, 0.035372, 
    0.035342, 0.035308, 0.035274, 0.035235, 0.035196, 0.035153, 0.035109, 
    0.035064, 0.035018, 0.034973, 0.034928, 0.034885, 0.034842, 0.034801, 
    0.034762, 0.034726, 0.034693, 0.034663, 0.034637, 0.034613, 0.034594, 
    0.034578, 0.034565, 0.034558, 0.034554, 0.034556, 0.034562, 0.034571, 
    0.034583, 0.034597, 0.034612, 0.034627, 0.034643, 0.034661, 0.034679, 
    0.034698, 0.034718, 0.034738, 0.034759, 0.034781, 0.034803, 0.034825, 
    0.034848, 0.03487, 0.034892, 0.034914, 0.034935, 0.030649, 0.030735, 
    0.030817, 0.030897, 0.030975, 0.03105, 0.031123, 0.031195, 0.031265, 
    0.031334, 0.031402, 0.03147, 0.031537, 0.031604, 0.031671, 0.031739, 
    0.031807, 0.031875, 0.031944, 0.032013, 0.032083, 0.032153, 0.032222, 
    0.032292, 0.032362, 0.03243, 0.032498, 0.032565, 0.03263, 0.032693, 
    0.032754, 0.032813, 0.03287, 0.032924, 0.032975, 0.033023, 0.033069, 
    0.033112, 0.033153, 0.03319, 0.033225, 0.033258, 0.033288, 0.033316, 
    0.033341, 0.033365, 0.033386, 0.033406, 0.033423, 0.033439, 0.033453, 
    0.033466, 0.033477, 0.033486, 0.033493, 0.033499, 0.033502, 0.033505, 
    0.033505, 0.033503, 0.0335, 0.033495, 0.033488, 0.033479, 0.033469, 
    0.033457, 0.033443, 0.033427, 0.033409, 0.033391, 0.03337, 0.033348, 
    0.033325, 0.0333, 0.033274, 0.033247, 0.033218, 0.033189, 0.033158, 
    0.033126, 0.033093, 0.033059, 0.033023, 0.032987, 0.032949, 0.03291, 
    0.03287, 0.032828, 0.032785, 0.032741, 0.032695, 0.032648, 0.032599, 
    0.03255, 0.032499, 0.032446, 0.032393, 0.032338, 0.032282, 0.032225, 
    0.032167, 0.032108, 0.032049, 0.031988, 0.031927, 0.031864, 0.031802, 
    0.031738, 0.031674, 0.031609, 0.031544, 0.031479, 0.031413, 0.031347, 
    0.03128, 0.031214, 0.031147, 0.03108, 0.031013, 0.030946, 0.03088, 
    0.030813, 0.030747, 0.03068, 0.030614, 0.030549, 0.030483, 0.030418, 
    0.030354, 0.030289, 0.030225, 0.030162, 0.030098, 0.030036, 0.029973, 
    0.029911, 0.029848, 0.029786, 0.029725, 0.029663, 0.029601, 0.02954, 
    0.029478, 0.029417, 0.029355, 0.029293, 0.029231, 0.029169, 0.029107, 
    0.029044, 0.028981, 0.028918, 0.028855, 0.028792, 0.028728, 0.028664, 
    0.028601, 0.028537, 0.028473, 0.02841, 0.028347, 0.028284, 0.028221, 
    0.028158, 0.028097, 0.028035, 0.027974, 0.027914, 0.027854, 0.027795, 
    0.027737, 0.027679, 0.027623, 0.027567, 0.027511, 0.027457, 0.027404, 
    0.027351, 0.0273, 0.027249, 0.027199, 0.02715, 0.027102, 0.027055, 
    0.027009, 0.026964, 0.026919, 0.026876, 0.026834, 0.026792, 0.026752, 
    0.026712, 0.026674, 0.026637, 0.0266, 0.026565, 0.026531, 0.026497, 
    0.026465, 0.026434, 0.026404, 0.026375, 0.026347, 0.02632, 0.026294, 
    0.026269, 0.026245, 0.026222, 0.026201, 0.02618, 0.026161, 0.026143, 
    0.026127, 0.026111, 0.026098, 0.026085, 0.026074, 0.026065, 0.026057, 
    0.026051, 0.026046, 0.026043, 0.026041, 0.02604, 0.026041, 0.026043, 
    0.026046, 0.02605, 0.026055, 0.026061, 0.026069, 0.026076, 0.026085, 
    0.026094, 0.026104, 0.026114, 0.026124, 0.026134, 0.026145, 0.026156, 
    0.026166, 0.026177, 0.026187, 0.026197, 0.026206, 0.026216, 0.026224, 
    0.026232, 0.02624, 0.026246, 0.026252, 0.026257, 0.026261, 0.026264, 
    0.026265, 0.026266, 0.026266, 0.026264, 0.026261, 0.026257, 0.026252, 
    0.026245, 0.026238, 0.026229, 0.026219, 0.026207, 0.026195, 0.026181, 
    0.026166, 0.02615, 0.026133, 0.026115, 0.026096, 0.026076, 0.026056, 
    0.026034, 0.026011, 0.025987, 0.025963, 0.025937, 0.02591, 0.025883, 
    0.025854, 0.025825, 0.025795, 0.025763, 0.025731, 0.025698, 0.025664, 
    0.025629, 0.025594, 0.025558, 0.025521, 0.025483, 0.025445, 0.025406, 
    0.025366, 0.025326, 0.025285, 0.025244, 0.025202, 0.025159, 0.025115, 
    0.025071, 0.025026, 0.02498, 0.024933, 0.024886, 0.024837, 0.024788, 
    0.024738, 0.024687, 0.024636, 0.024583, 0.02453, 0.024477, 0.024423, 
    0.024368, 0.024313, 0.024258, 0.024202, 0.024147, 0.024092, 0.024036, 
    0.023981, 0.023926, 0.023872, 0.023819, 0.023766, 0.023714, 0.023663, 
    0.023613, 0.023565, 0.023518, 0.023473, 0.02343, 0.023389, 0.02335, 
    0.023314, 0.023279, 0.023248, 0.023219, 0.023192, 0.023168, 0.023146, 
    0.023126, 0.023109, 0.023093, 0.02308, 0.023068, 0.023058, 0.02305, 
    0.023043, 0.023037, 0.023033, 0.02303, 0.023028, 0.023027, 0.023027, 
    0.023028, 0.02303, 0.023032, 0.023035, 0.023038, 0.023041, 0.023045, 
    0.023049, 0.023053, 0.023058, 0.023062, 0.023066, 0.02307, 0.023074, 
    0.023078, 0.023081, 0.023084, 0.023086, 0.023088, 0.02309, 0.023091, 
    0.023091, 0.02309, 0.023089, 0.023087, 0.023084, 0.023079, 0.023074, 
    0.023068, 0.023061, 0.023053, 0.023043, 0.023032, 0.02302, 0.023006, 
    0.022991, 0.022975, 0.022958, 0.022939, 0.022919, 0.022898, 0.022876, 
    0.022852, 0.022827, 0.022801, 0.022774, 0.022746, 0.022716, 0.022685, 
    0.022653, 0.02262, 0.022585, 0.02255, 0.022513, 0.022474, 0.022435, 
    0.022395, 0.022354, 0.022312, 0.022269, 0.022225, 0.02218, 0.022135, 
    0.02209, 0.022044, 0.021998, 0.021951, 0.021905, 0.021858, 0.021811, 
    0.021765, 0.021718, 0.021672, 0.021625, 0.021579, 0.021534, 0.021488, 
    0.021443, 0.021398, 0.021353, 0.021309, 0.021265, 0.021222, 0.021179, 
    0.021137, 0.021095, 0.021054, 0.021014, 0.020975, 0.020936, 0.020898, 
    0.020862, 0.020826, 0.020792, 0.020758, 0.020726, 0.020696, 0.020666, 
    0.020637, 0.02061, 0.020584, 0.020558, 0.020534, 0.02051, 0.020487, 
    0.020465, 0.020444, 0.020424, 0.020404, 0.020385, 0.020367, 0.020349, 
    0.020332, 0.020315, 0.020299, 0.020284, 0.020269, 0.020254, 0.020239, 
    0.020225, 0.020211, 0.020198, 0.020184, 0.02017, 0.020157, 0.020143, 
    0.02013, 0.020116, 0.020102, 0.020088, 0.020073, 0.020058, 0.020043, 
    0.020027, 0.020011, 0.019994, 0.019977, 0.019959, 0.01994, 0.019921, 
    0.019902, 0.019882, 0.019862, 0.019842, 0.019822, 0.019801, 0.01978, 
    0.019758, 0.019737, 0.019715, 0.019693, 0.019671, 0.019648, 0.019625, 
    0.019602, 0.019579, 0.019555, 0.019531, 0.019506, 0.019482, 0.019456, 
    0.019431, 0.019405, 0.019379, 0.019352, 0.019325, 0.019298, 0.01927, 
    0.019243, 0.019215, 0.019187, 0.019159, 0.019131, 0.019103, 0.019076, 
    0.019048, 0.019021, 0.018994, 0.018968, 0.018942, 0.018916, 0.018892, 
    0.018868, 0.018844, 0.018822, 0.018801, 0.01878, 0.01876, 0.018742, 
    0.018724, 0.018708, 0.018692, 0.018677, 0.018663, 0.018649, 0.018636, 
    0.018624, 0.018613, 0.018602, 0.018591, 0.018581, 0.018571, 0.018562, 
    0.018553, 0.018545, 0.018536, 0.018528, 0.01852, 0.018512, 0.018504, 
    0.018496, 0.018488, 0.018481, 0.018473, 0.018465, 0.018457, 0.018448, 
    0.01844, 0.018431, 0.018422, 0.018413, 0.018403, 0.018393, 0.018383, 
    0.018372, 0.01836, 0.018348, 0.018336, 0.018322, 0.018308, 0.018293, 
    0.018278, 0.018262, 0.018245, 0.018227, 0.018209, 0.01819, 0.01817, 
    0.01815, 0.018129, 0.018107, 0.018085, 0.018062, 0.018038, 0.018014, 
    0.017989, 0.017964, 0.017938, 0.017912, 0.017885, 0.017858, 0.01783, 
    0.017802, 0.017774, 0.017745, 0.017717, 0.017688, 0.017659, 0.01763, 
    0.017601, 0.017573, 0.017544, 0.017516, 0.017488, 0.01746, 0.017433, 
    0.017407, 0.017381, 0.017355, 0.01733, 0.017306, 0.017282, 0.017259, 
    0.017237, 0.017216, 0.017195, 0.017175, 0.017156, 0.017137, 0.017119, 
    0.017101, 0.017084, 0.017067, 0.017051, 0.017035, 0.017019, 0.017003, 
    0.016988, 0.016973, 0.016959, 0.016944, 0.016929, 0.016915, 0.0169, 
    0.016886, 0.016871, 0.016857, 0.016842, 0.016827, 0.016812, 0.016796, 
    0.016781, 0.016765, 0.016748, 0.016732, 0.016715, 0.016697, 0.01668, 
    0.016661, 0.016643, 0.016623, 0.016604, 0.016583, 0.016562, 0.016541, 
    0.016519, 0.016495, 0.016472, 0.016447, 0.016422, 0.016396, 0.01637, 
    0.016342, 0.016314, 0.016286, 0.016257, 0.016227, 0.016197, 0.016166, 
    0.016135, 0.016104, 0.016072, 0.016039, 0.016007, 0.015974, 0.015941, 
    0.015908, 0.015875, 0.015842, 0.015809, 0.015776, 0.015744, 0.015712, 
    0.015681, 0.01565, 0.01562, 0.015591, 0.015563, 0.015536, 0.015511, 
    0.015486, 0.015463, 0.015442, 0.015421, 0.015402, 0.015385, 0.015368, 
    0.015352, 0.015338, 0.015324, 0.015311, 0.015299, 0.015287, 0.015276, 
    0.015266, 0.015256, 0.015247, 0.015238, 0.015229, 0.01522, 0.015212, 
    0.015203, 0.015195, 0.015186, 0.015178, 0.015169, 0.01516, 0.01515, 
    0.01514, 0.01513, 0.015119, 0.015108, 0.015096, 0.015083, 0.01507, 
    0.015056, 0.01504, 0.015024, 0.015008, 0.01499, 0.014972, 0.014953, 
    0.014934, 0.014913, 0.014892, 0.014871, 0.014849, 0.014826, 0.014803, 
    0.014779, 0.014755, 0.01473, 0.014705, 0.01468, 0.014654, 0.014628, 
    0.014601, 0.014574, 0.014547, 0.01452, 0.014492, 0.014464, 0.014436, 
    0.014408, 0.01438, 0.014351, 0.014323, 0.014295, 0.014266, 0.014237, 
    0.014209, 0.01418, 0.014152, 0.014123, 0.014095, 0.014066, 0.014038, 
    0.014009, 0.013981, 0.013953, 0.013924, 0.013896, 0.013868, 0.01384, 
    0.013811, 0.013783, 0.013755, 0.013727, 0.013698, 0.01367, 0.013642, 
    0.013614, 0.013585, 0.013557, 0.013529, 0.013501, 0.013473, 0.013445, 
    0.013418, 0.01339, 0.013362, 0.013335, 0.013307, 0.01328, 0.013253, 
    0.013225, 0.013198, 0.013171, 0.013144, 0.013117, 0.013091, 0.013064, 
    0.013037, 0.01301, 0.012984, 0.012957, 0.012931, 0.012904, 0.012878, 
    0.012851, 0.012825, 0.012798, 0.012772, 0.012745, 0.012718, 0.012692, 
    0.012665, 0.012638, 0.012611, 0.012584, 0.012557, 0.01253, 0.012502, 
    0.012475, 0.012447, 0.01242, 0.012392, 0.012364, 0.012336, 0.012308, 
    0.01228, 0.012251, 0.012223, 0.012194, 0.012165, 0.012137, 0.012108, 
    0.012079, 0.01205, 0.012021, 0.011991, 0.011962, 0.011933, 0.011903, 
    0.011874, 0.011844, 0.011814, 0.011785, 0.011755, 0.011725, 0.011695, 
    0.011665, 0.011635, 0.011605, 0.011574, 0.011544, 0.011514, 0.011483, 
    0.011453, 0.011422, 0.011391, 0.011361, 0.01133, 0.0113, 0.011269, 
    0.011238, 0.011208, 0.011177, 0.011147, 0.011116, 0.011086, 0.011055, 
    0.011025, 0.010995, 0.010965, 0.010935, 0.010905, 0.010875, 0.010845, 
    0.010815, 0.010785, 0.010755, 0.010725, 0.010695, 0.010665, 0.010635, 
    0.010604, 0.010574, 0.010544, 0.010514, 0.010483, 0.010453, 0.010422, 
    0.010391, 0.01036, 0.010329, 0.010298, 0.010267, 0.010235, 0.010204, 
    0.010172, 0.01014, 0.010107, 0.010075, 0.010042, 0.010009, 0.0099763, 
    0.009943, 0.0099095, 0.0098759, 0.009842, 0.009808, 0.0097737, 0.0097393, 
    0.0097047, 0.0096699, 0.009635, 0.0095999, 0.0095647, 0.0095294, 
    0.0094939, 0.0094584, 0.0094229, 0.0093873, 0.0093517, 0.0093161, 
    0.0092805, 0.009245, 0.0092094, 0.009174, 0.0091386, 0.0091033, 0.009068, 
    0.0090328, 0.0089977, 0.0089626, 0.0089276, 0.0088926, 0.0088577, 
    0.0088228, 0.0087879, 0.0087529, 0.008718, 0.008683, 0.008648, 0.008613, 
    0.0085779, 0.0085428, 0.0085076, 0.0084724, 0.0084372, 0.0084019, 
    0.0083667, 0.0083314, 0.0082961, 0.0082609, 0.0082256, 0.0081904, 
    0.0081552, 0.00812, 0.0080849, 0.0080498, 0.0080148, 0.0079798, 
    0.0079449, 0.0079101, 0.0078753, 0.0078407, 0.0078061, 0.0077716, 
    0.0077372, 0.0077029, 0.0076687, 0.0076346, 0.0076007, 0.0075668, 
    0.0075331, 0.0074995, 0.0074659, 0.0074325, 0.0073992, 0.007366, 
    0.0073329, 0.0072999, 0.007267, 0.0072342, 0.0072015, 0.0071688, 
    0.0071362, 0.0071037, 0.0070712, 0.0070388, 0.0070065, 0.0069742, 
    0.0069419, 0.0069098, 0.0068777, 0.0068457, 0.0068137, 0.0067818, 
    0.00675, 0.0067183, 0.0066867, 0.0066552, 0.0066238, 0.0065925, 
    0.0065613, 0.0065302, 0.0064992, 0.0064683, 0.0064375, 0.0064069, 
    0.0063764, 0.006346, 0.0063157, 0.0062855, 0.0062555, 0.0062257, 
    0.006196, 0.0061664, 0.0061369, 0.0061076, 0.0060785, 0.0060494, 
    0.0060205, 0.0059918, 0.0059631, 0.0059346, 0.0059061, 0.0058778, 
    0.0058495, 0.0058213, 0.0057932, 0.0057652, 0.0057373, 0.0057094, 
    0.0056816, 0.0056538, 0.0056261, 0.0055985, 0.005571, 0.0055435, 
    0.0055161, 0.0054888, 0.0054616, 0.0054344, 0.0054074, 0.0053804, 
    0.0053535, 0.0053266, 0.0052999, 0.0052732, 0.0052466, 0.0052201, 
    0.0051937, 0.0051673, 0.005141, 0.0051148, 0.0050887, 0.0050626, 
    0.0050366, 0.0050107, 0.0049849, 0.0049592, 0.0049335, 0.0049079, 
    0.0048825, 0.0048571, 0.0048318, 0.0048067, 0.0047816, 0.0047566, 
    0.0047318, 0.004707, 0.0046824, 0.0046578, 0.0046334, 0.0046091, 
    0.0045848, 0.0045607, 0.0045367, 0.0045127, 0.0044889, 0.0044651, 
    0.0044415, 0.0044179, 0.0043945, 0.0043711, 0.0043478, 0.0043247, 
    0.0043016, 0.0042786, 0.0042557, 0.004233, 0.0042103, 0.0041877, 
    0.0041653, 0.0041429, 0.0041207, 0.0040985, 0.0040765, 0.0040546, 
    0.0040328, 0.0040111, 0.0039895, 0.0039681, 0.0039467, 0.0039255, 
    0.0039043, 0.0038833, 0.0038624, 0.0038416, 0.0038209, 0.0038003, 
    0.0037799, 0.0037595, 0.0037392, 0.0037191, 0.0036991, 0.0036792, 
    0.0036593, 0.0036396, 0.00362, 0.0036005, 0.0035811, 0.0035618, 
    0.0035426, 0.0035235, 0.0035044, 0.0034855, 0.0034666, 0.0034478, 
    0.0034291, 0.0034105, 0.003392, 0.0033735, 0.0033551, 0.0033368, 
    0.0033186, 0.0033005, 0.0032825, 0.0032645, 0.0032466, 0.0032289, 
    0.0032112, 0.0031936, 0.0031761, 0.0031587, 0.0031414, 0.0031242, 
    0.0031071, 0.0030901, 0.0030732, 0.0030564, 0.0030398, 0.0030232, 
    0.0030067, 0.0029903, 0.0029741, 0.0029579, 0.0029419, 0.002926, 
    0.0029102, 0.0028944, 0.0028789, 0.0028634, 0.002848, 0.0028327, 
    0.0028176, 0.0028025, 0.0027875, 0.0027727, 0.0027579, 0.0027432, 
    0.0027286, 0.0027141, 0.0026997, 0.0026853, 0.002671, 0.0026567, 
    0.0026425, 0.0026284, 0.0026143, 0.0026003, 0.0025863, 0.0025724, 
    0.0025586, 0.0025448, 0.0025311, 0.0025174, 0.0025039, 0.0024904, 
    0.002477, 0.0024637, 0.0024505, 0.0024374, 0.0024244, 0.0024116, 
    0.0023988, 0.0023862, 0.0023737, 0.0023614, 0.0023491, 0.002337, 
    0.002325, 0.0023132, 0.0023014, 0.0022898, 0.0022782, 0.0022668, 
    0.0022554, 0.0022441, 0.0022329, 0.0022218, 0.0022107, 0.0021997, 
    0.0021888, 0.0021778, 0.0021669, 0.0021561, 0.0021452, 0.0021344, 
    0.0021236, 0.0021129, 0.0021021, 0.0020914, 0.0020807, 0.0020701, 
    0.0020594, 0.0020488, 0.0020382, 0.0020277, 0.0020171, 0.0020067, 
    0.0019963, 0.0019859, 0.0019756, 0.0019653, 0.0019551, 0.001945, 
    0.0019349, 0.0019249, 0.001915, 0.0019051, 0.0018953, 0.0018857, 
    0.0018761, 0.0018665, 0.0018571, 0.0018478, 0.0018385, 0.0018293, 
    0.0018202, 0.0018113, 0.0018024, 0.0017935, 0.0017848, 0.0017761, 
    0.0017676, 0.001759, 0.0017506, 0.0017422, 0.0017339, 0.0017257, 
    0.0017175, 0.0017094, 0.0017013, 0.0016933, 0.0016854, 0.0016775, 
    0.0016697, 0.0016619, 0.0016542, 0.0016465, 0.0016389, 0.0016313, 
    0.0016238, 0.0016164, 0.001609, 0.0016017, 0.0015945, 0.0015874, 
    0.0015803, 0.0015733, 0.0015663, 0.0015594, 0.0015527, 0.0015459, 
    0.0015393, 0.0015328, 0.0015263, 0.0015199, 0.0015136, 0.0015073, 
    0.0015011, 0.001495, 0.0014889, 0.0014829, 0.001477, 0.0014711, 
    0.0014653, 0.0014595, 0.0014537, 0.001448, 0.0014423, 0.0014367, 
    0.0014311, 0.0014255, 0.00142, 0.0014145, 0.001409, 0.0014036, 0.0013981, 
    0.0013927, 0.0013873, 0.0013819, 0.0013765, 0.0013712, 0.0013658, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 refrac_qual =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100 ;

 dry_temp =
  267.89, 267.63, 267.36, 267.09, 266.81, 266.53, 266.26, 265.99, 265.72, 
    265.46, 265.2, 264.95, 264.71, 264.49, 264.27, 264.07, 263.88, 263.71, 
    263.55, 263.4, 263.26, 263.14, 263.03, 262.93, 262.84, 262.74, 262.65, 
    262.57, 262.49, 262.42, 262.34, 262.27, 262.21, 262.14, 262.09, 262.04, 
    262, 261.96, 261.93, 261.91, 261.89, 261.87, 261.86, 261.85, 261.85, 
    261.84, 261.84, 261.83, 261.82, 261.82, 261.81, 261.8, 261.79, 261.77, 
    261.76, 261.74, 261.73, 261.71, 261.68, 261.66, 261.64, 261.62, 261.61, 
    261.6, 261.59, 261.58, 261.57, 261.55, 261.54, 261.53, 261.51, 261.5, 
    261.48, 261.46, 261.44, 261.41, 261.39, 261.36, 261.33, 261.3, 261.26, 
    261.23, 261.19, 261.15, 261.12, 261.08, 261.05, 261.02, 260.99, 260.97, 
    260.94, 260.92, 260.89, 260.87, 260.85, 260.84, 260.82, 260.81, 260.79, 
    260.78, 260.77, 260.76, 260.75, 260.74, 260.73, 260.73, 260.72, 260.72, 
    260.71, 260.71, 260.7, 260.7, 260.69, 260.69, 260.69, 260.69, 260.69, 
    260.69, 260.68, 260.68, 260.68, 260.67, 260.66, 260.65, 260.64, 260.63, 
    260.62, 260.6, 260.59, 260.57, 260.55, 260.54, 260.52, 260.51, 260.49, 
    260.47, 260.46, 260.44, 260.43, 260.42, 260.4, 260.39, 260.38, 260.37, 
    260.36, 260.34, 260.33, 260.32, 260.31, 260.29, 260.28, 260.27, 260.26, 
    260.25, 260.23, 260.22, 260.22, 260.21, 260.2, 260.2, 260.19, 260.2, 
    260.2, 260.21, 260.22, 260.23, 260.25, 260.27, 260.29, 260.31, 260.34, 
    260.36, 260.4, 260.43, 260.47, 260.51, 260.55, 260.59, 260.64, 260.69, 
    260.74, 260.8, 260.87, 260.94, 261.02, 261.1, 261.2, 261.31, 261.43, 
    261.56, 261.7, 261.86, 262.02, 262.19, 262.36, 262.53, 262.71, 262.88, 
    263.05, 263.21, 263.38, 263.53, 263.69, 263.85, 264.01, 264.17, 264.34, 
    264.5, 264.67, 264.84, 265.01, 265.17, 265.34, 265.51, 265.68, 265.84, 
    265.99, 266.14, 266.28, 266.42, 266.55, 266.68, 266.8, 266.92, 267.02, 
    267.11, 267.19, 267.26, 267.31, 267.35, 267.38, 267.41, 267.43, 267.45, 
    267.48, 267.5, 267.53, 267.57, 267.61, 267.65, 267.7, 267.75, 267.79, 
    267.83, 267.87, 267.9, 267.93, 267.95, 267.98, 268, 268.01, 268.01, 
    268.01, 268, 268, 268.01, 268.02, 268.02, 268.02, 268.02, 268.02, 268.01, 
    267.99, 267.96, 267.94, 267.92, 267.89, 267.86, 267.82, 267.78, 267.74, 
    267.7, 267.65, 267.59, 267.53, 267.47, 267.41, 267.33, 267.25, 267.17, 
    267.09, 267.01, 266.93, 266.84, 266.75, 266.66, 266.57, 266.48, 266.4, 
    266.31, 266.23, 266.16, 266.08, 266, 265.92, 265.84, 265.77, 265.69, 
    265.62, 265.54, 265.48, 265.43, 265.37, 265.32, 265.28, 265.23, 265.19, 
    265.15, 265.11, 265.07, 265.03, 264.99, 264.96, 264.92, 264.88, 264.84, 
    264.79, 264.75, 264.71, 264.66, 264.62, 264.57, 264.53, 264.49, 264.46, 
    264.42, 264.39, 264.36, 264.33, 264.29, 264.26, 264.22, 264.18, 264.13, 
    264.08, 264.03, 263.98, 263.92, 263.85, 263.78, 263.7, 263.62, 263.54, 
    263.45, 263.37, 263.28, 263.19, 263.11, 263.03, 262.95, 262.87, 262.79, 
    262.72, 262.64, 262.58, 262.51, 262.44, 262.38, 262.32, 262.26, 262.19, 
    262.13, 262.06, 261.99, 261.92, 261.85, 261.78, 261.71, 261.64, 261.58, 
    261.52, 261.46, 261.4, 261.35, 261.3, 261.25, 261.21, 261.17, 261.14, 
    261.11, 261.08, 261.05, 261.02, 260.99, 260.97, 260.94, 260.91, 260.89, 
    260.86, 260.84, 260.81, 260.79, 260.76, 260.74, 260.72, 260.7, 260.68, 
    260.66, 260.65, 260.63, 260.61, 260.59, 260.57, 260.55, 260.53, 260.5, 
    260.48, 260.45, 260.43, 260.4, 260.37, 260.34, 260.31, 260.28, 260.25, 
    260.22, 260.19, 260.16, 260.13, 260.1, 260.07, 260.04, 260.01, 259.98, 
    259.95, 259.92, 259.89, 259.86, 259.82, 259.79, 259.75, 259.72, 259.68, 
    259.65, 259.61, 259.57, 259.54, 259.5, 259.46, 259.43, 259.4, 259.37, 
    259.34, 259.31, 259.28, 259.25, 259.23, 259.2, 259.17, 259.14, 259.11, 
    259.08, 259.05, 259.02, 258.99, 258.95, 258.92, 258.89, 258.86, 258.82, 
    258.79, 258.75, 258.72, 258.69, 258.66, 258.63, 258.6, 258.57, 258.53, 
    258.5, 258.47, 258.44, 258.4, 258.37, 258.33, 258.3, 258.26, 258.22, 
    258.17, 258.13, 258.08, 258.04, 258, 257.96, 257.92, 257.88, 257.84, 
    257.8, 257.77, 257.74, 257.7, 257.68, 257.65, 257.62, 257.59, 257.56, 
    257.54, 257.51, 257.49, 257.46, 257.44, 257.41, 257.38, 257.35, 257.32, 
    257.3, 257.27, 257.24, 257.22, 257.19, 257.17, 257.14, 257.12, 257.09, 
    257.07, 257.05, 257.04, 257.02, 257, 256.98, 256.96, 256.94, 256.93, 
    256.91, 256.89, 256.87, 256.85, 256.83, 256.81, 256.79, 256.77, 256.75, 
    256.73, 256.71, 256.69, 256.67, 256.65, 256.63, 256.61, 256.6, 256.58, 
    256.56, 256.54, 256.52, 256.51, 256.49, 256.47, 256.45, 256.43, 256.41, 
    256.39, 256.37, 256.35, 256.33, 256.31, 256.29, 256.27, 256.25, 256.23, 
    256.21, 256.18, 256.16, 256.14, 256.12, 256.09, 256.07, 256.04, 256.02, 
    256, 255.97, 255.95, 255.93, 255.91, 255.89, 255.87, 255.85, 255.83, 
    255.81, 255.79, 255.78, 255.77, 255.75, 255.74, 255.73, 255.72, 255.71, 
    255.7, 255.69, 255.68, 255.67, 255.66, 255.65, 255.64, 255.63, 255.62, 
    255.61, 255.6, 255.59, 255.58, 255.58, 255.57, 255.56, 255.55, 255.54, 
    255.54, 255.53, 255.52, 255.52, 255.51, 255.5, 255.49, 255.48, 255.46, 
    255.45, 255.43, 255.42, 255.4, 255.38, 255.35, 255.33, 255.31, 255.29, 
    255.27, 255.24, 255.22, 255.19, 255.17, 255.14, 255.12, 255.1, 255.08, 
    255.05, 255.03, 255.01, 254.99, 254.97, 254.95, 254.93, 254.91, 254.89, 
    254.87, 254.85, 254.83, 254.81, 254.79, 254.76, 254.74, 254.71, 254.68, 
    254.66, 254.63, 254.6, 254.58, 254.55, 254.52, 254.49, 254.47, 254.44, 
    254.41, 254.38, 254.35, 254.32, 254.29, 254.27, 254.24, 254.21, 254.18, 
    254.15, 254.13, 254.1, 254.07, 254.04, 254.01, 253.98, 253.95, 253.91, 
    253.88, 253.84, 253.81, 253.77, 253.73, 253.7, 253.66, 253.63, 253.6, 
    253.57, 253.54, 253.51, 253.48, 253.45, 253.43, 253.41, 253.39, 253.38, 
    253.36, 253.35, 253.34, 253.33, 253.32, 253.31, 253.3, 253.29, 253.29, 
    253.28, 253.28, 253.27, 253.27, 253.26, 253.25, 253.24, 253.23, 253.22, 
    253.21, 253.21, 253.2, 253.19, 253.18, 253.17, 253.16, 253.15, 253.15, 
    253.14, 253.13, 253.12, 253.11, 253.1, 253.09, 253.07, 253.06, 253.05, 
    253.03, 253.01, 253, 252.98, 252.96, 252.94, 252.92, 252.9, 252.88, 
    252.86, 252.84, 252.81, 252.79, 252.76, 252.73, 252.71, 252.68, 252.66, 
    252.63, 252.61, 252.58, 252.55, 252.53, 252.5, 252.48, 252.45, 252.43, 
    252.4, 252.37, 252.35, 252.32, 252.29, 252.26, 252.23, 252.2, 252.17, 
    252.14, 252.11, 252.09, 252.06, 252.04, 252.02, 252.01, 252, 251.99, 
    251.99, 251.99, 251.99, 252, 252.01, 252.02, 252.03, 252.05, 252.07, 
    252.09, 252.11, 252.14, 252.17, 252.2, 252.24, 252.28, 252.32, 252.36, 
    252.41, 252.46, 252.52, 252.57, 252.63, 252.7, 252.76, 252.84, 252.91, 
    252.99, 253.07, 253.15, 253.24, 253.33, 253.42, 253.52, 253.62, 253.71, 
    253.81, 253.9, 254, 254.1, 254.2, 254.3, 254.4, 254.5, 254.6, 254.7, 
    254.8, 254.9, 255.01, 255.11, 255.21, 255.31, 255.41, 255.51, 255.6, 
    255.7, 255.79, 255.88, 255.97, 256.06, 256.15, 256.23, 256.31, 256.38, 
    256.46, 256.53, 256.59, 256.65, 256.71, 256.77, 256.81, 256.86, 256.9, 
    256.93, 256.96, 256.99, 257.01, 257.03, 257.04, 257.05, 257.06, 257.06, 
    257.07, 257.07, 257.07, 257.07, 257.07, 257.06, 257.05, 257.04, 257.03, 
    257.01, 257, 256.99, 256.97, 256.95, 256.94, 256.92, 256.91, 256.89, 
    256.88, 256.87, 256.85, 256.84, 256.83, 256.82, 256.81, 256.8, 256.79, 
    256.78, 256.77, 256.76, 256.76, 256.75, 256.74, 256.73, 256.73, 256.72, 
    256.71, 256.7, 256.69, 256.68, 256.67, 256.66, 256.65, 256.64, 256.63, 
    256.62, 256.61, 256.59, 256.58, 256.57, 256.56, 256.55, 256.53, 256.52, 
    256.51, 256.5, 256.48, 256.47, 256.46, 256.44, 256.43, 256.41, 256.4, 
    256.38, 256.36, 256.34, 256.32, 256.3, 256.28, 256.25, 256.23, 256.2, 
    256.18, 256.15, 256.12, 256.09, 256.07, 256.04, 256.01, 255.98, 255.95, 
    255.92, 255.89, 255.86, 255.83, 255.8, 255.77, 255.74, 255.71, 255.68, 
    255.65, 255.62, 255.59, 255.56, 255.53, 255.5, 255.46, 255.43, 255.4, 
    255.36, 255.33, 255.3, 255.26, 255.23, 255.2, 255.17, 255.14, 255.11, 
    255.08, 255.05, 255.02, 254.99, 254.96, 254.93, 254.89, 254.86, 254.83, 
    254.8, 254.76, 254.73, 254.69, 254.66, 254.62, 254.59, 254.55, 254.52, 
    254.48, 254.45, 254.42, 254.38, 254.35, 254.32, 254.29, 254.26, 254.23, 
    254.19, 254.16, 254.13, 254.1, 254.07, 254.04, 254.01, 253.98, 253.95, 
    253.92, 253.89, 253.87, 253.84, 253.81, 253.78, 253.76, 253.73, 253.71, 
    253.68, 253.66, 253.64, 253.62, 253.6, 253.58, 253.56, 253.54, 253.53, 
    253.51, 253.49, 253.48, 253.46, 253.45, 253.44, 253.42, 253.41, 253.39, 
    253.37, 253.36, 253.34, 253.33, 253.31, 253.29, 253.27, 253.26, 253.24, 
    253.22, 253.2, 253.18, 253.16, 253.14, 253.12, 253.1, 253.08, 253.07, 
    253.05, 253.03, 253.01, 252.99, 252.97, 252.95, 252.93, 252.91, 252.89, 
    252.87, 252.84, 252.82, 252.8, 252.77, 252.74, 252.71, 252.68, 252.66, 
    252.63, 252.6, 252.57, 252.54, 252.51, 252.48, 252.45, 252.43, 252.4, 
    252.37, 252.35, 252.32, 252.29, 252.27, 252.24, 252.21, 252.19, 252.16, 
    252.13, 252.1, 252.07, 252.04, 252.01, 251.99, 251.96, 251.93, 251.9, 
    251.87, 251.84, 251.82, 251.79, 251.76, 251.74, 251.71, 251.68, 251.66, 
    251.64, 251.61, 251.59, 251.56, 251.54, 251.52, 251.5, 251.47, 251.45, 
    251.43, 251.41, 251.39, 251.37, 251.35, 251.34, 251.32, 251.3, 251.29, 
    251.27, 251.25, 251.23, 251.22, 251.2, 251.19, 251.17, 251.15, 251.14, 
    251.12, 251.11, 251.09, 251.07, 251.06, 251.04, 251.02, 251, 250.99, 
    250.97, 250.95, 250.93, 250.92, 250.9, 250.88, 250.86, 250.84, 250.82, 
    250.8, 250.77, 250.75, 250.73, 250.7, 250.68, 250.65, 250.62, 250.59, 
    250.56, 250.53, 250.5, 250.47, 250.45, 250.42, 250.39, 250.36, 250.33, 
    250.3, 250.27, 250.24, 250.21, 250.17, 250.14, 250.11, 250.08, 250.05, 
    250.02, 249.98, 249.95, 249.92, 249.88, 249.85, 249.82, 249.79, 249.76, 
    249.72, 249.69, 249.66, 249.63, 249.6, 249.57, 249.54, 249.5, 249.48, 
    249.45, 249.42, 249.39, 249.37, 249.34, 249.32, 249.3, 249.27, 249.25, 
    249.22, 249.2, 249.17, 249.15, 249.12, 249.1, 249.08, 249.05, 249.03, 
    249, 248.98, 248.95, 248.93, 248.91, 248.88, 248.86, 248.84, 248.81, 
    248.79, 248.77, 248.74, 248.72, 248.7, 248.68, 248.66, 248.64, 248.62, 
    248.6, 248.58, 248.56, 248.54, 248.52, 248.5, 248.48, 248.45, 248.43, 
    248.41, 248.39, 248.36, 248.34, 248.31, 248.29, 248.26, 248.24, 248.21, 
    248.19, 248.16, 248.14, 248.11, 248.09, 248.06, 248.04, 248.01, 247.98, 
    247.96, 247.93, 247.91, 247.88, 247.85, 247.83, 247.8, 247.77, 247.74, 
    247.71, 247.68, 247.65, 247.61, 247.58, 247.55, 247.51, 247.48, 247.44, 
    247.41, 247.38, 247.34, 247.31, 247.28, 247.25, 247.22, 247.19, 247.16, 
    247.13, 247.1, 247.08, 247.05, 247.02, 246.99, 246.97, 246.94, 246.91, 
    246.89, 246.87, 246.84, 246.82, 246.8, 246.78, 246.76, 246.74, 246.71, 
    246.69, 246.67, 246.65, 246.63, 246.62, 246.6, 246.58, 246.56, 246.54, 
    246.52, 246.5, 246.48, 246.46, 246.44, 246.42, 246.41, 246.39, 246.37, 
    246.35, 246.33, 246.31, 246.3, 246.28, 246.26, 246.24, 246.23, 246.21, 
    246.19, 246.17, 246.15, 246.13, 246.11, 246.09, 246.07, 246.04, 246.02, 
    246, 245.98, 245.96, 245.94, 245.92, 245.9, 245.88, 245.87, 245.85, 
    245.83, 245.81, 245.79, 245.77, 245.75, 245.73, 245.71, 245.69, 245.67, 
    245.64, 245.62, 245.6, 245.58, 245.56, 245.54, 245.51, 245.49, 245.47, 
    245.45, 245.43, 245.4, 245.38, 245.36, 245.34, 245.32, 245.3, 245.28, 
    245.26, 245.24, 245.22, 245.2, 245.18, 245.16, 245.14, 245.12, 245.1, 
    245.08, 245.06, 245.04, 245.02, 245, 244.98, 244.96, 244.94, 244.92, 
    244.9, 244.89, 244.87, 244.85, 244.84, 244.82, 244.8, 244.79, 244.77, 
    244.75, 244.73, 244.72, 244.7, 244.68, 244.67, 244.65, 244.64, 244.63, 
    244.61, 244.6, 244.58, 244.56, 244.55, 244.53, 244.51, 244.49, 244.47, 
    244.45, 244.43, 244.41, 244.39, 244.37, 244.35, 244.33, 244.31, 244.29, 
    244.27, 244.25, 244.22, 244.2, 244.18, 244.15, 244.13, 244.1, 244.08, 
    244.05, 244.02, 243.99, 243.96, 243.94, 243.91, 243.88, 243.85, 243.82, 
    243.79, 243.75, 243.72, 243.69, 243.66, 243.63, 243.6, 243.57, 243.54, 
    243.51, 243.48, 243.45, 243.42, 243.39, 243.36, 243.33, 243.3, 243.27, 
    243.24, 243.21, 243.18, 243.15, 243.12, 243.09, 243.07, 243.04, 243.01, 
    242.98, 242.96, 242.93, 242.9, 242.87, 242.85, 242.82, 242.8, 242.77, 
    242.75, 242.72, 242.7, 242.67, 242.64, 242.62, 242.59, 242.57, 242.54, 
    242.51, 242.49, 242.46, 242.43, 242.41, 242.38, 242.35, 242.33, 242.3, 
    242.27, 242.25, 242.22, 242.19, 242.17, 242.14, 242.11, 242.09, 242.06, 
    242.03, 242, 241.97, 241.95, 241.92, 241.89, 241.86, 241.83, 241.81, 
    241.78, 241.75, 241.72, 241.7, 241.67, 241.64, 241.62, 241.59, 241.57, 
    241.54, 241.52, 241.49, 241.47, 241.44, 241.42, 241.4, 241.37, 241.35, 
    241.33, 241.3, 241.28, 241.26, 241.24, 241.21, 241.19, 241.17, 241.14, 
    241.12, 241.1, 241.07, 241.05, 241.03, 241.01, 240.98, 240.96, 240.94, 
    240.91, 240.89, 240.86, 240.83, 240.81, 240.78, 240.75, 240.73, 240.7, 
    240.67, 240.64, 240.62, 240.59, 240.56, 240.53, 240.51, 240.48, 240.45, 
    240.42, 240.4, 240.37, 240.34, 240.32, 240.29, 240.26, 240.23, 240.2, 
    240.17, 240.14, 240.11, 240.08, 240.05, 240.02, 239.99, 239.96, 239.93, 
    239.9, 239.87, 239.85, 239.82, 239.79, 239.76, 239.74, 239.71, 239.68, 
    239.65, 239.63, 239.6, 239.57, 239.54, 239.52, 239.49, 239.46, 239.43, 
    239.4, 239.37, 239.34, 239.31, 239.28, 239.25, 239.22, 239.19, 239.16, 
    239.14, 239.11, 239.08, 239.05, 239.02, 238.99, 238.96, 238.94, 238.91, 
    238.88, 238.86, 238.83, 238.8, 238.77, 238.75, 238.72, 238.69, 238.66, 
    238.64, 238.61, 238.58, 238.56, 238.53, 238.5, 238.47, 238.44, 238.41, 
    238.38, 238.36, 238.33, 238.3, 238.27, 238.25, 238.22, 238.19, 238.16, 
    238.13, 238.11, 238.08, 238.05, 238.03, 238, 237.98, 237.95, 237.92, 
    237.9, 237.88, 237.85, 237.83, 237.81, 237.78, 237.76, 237.74, 237.72, 
    237.7, 237.67, 237.65, 237.63, 237.61, 237.59, 237.57, 237.55, 237.53, 
    237.51, 237.49, 237.47, 237.45, 237.43, 237.41, 237.39, 237.37, 237.35, 
    237.33, 237.31, 237.29, 237.27, 237.26, 237.24, 237.22, 237.2, 237.18, 
    237.16, 237.15, 237.13, 237.11, 237.09, 237.07, 237.05, 237.03, 237.01, 
    236.99, 236.96, 236.94, 236.92, 236.9, 236.87, 236.85, 236.82, 236.8, 
    236.77, 236.75, 236.73, 236.7, 236.68, 236.66, 236.63, 236.61, 236.59, 
    236.56, 236.54, 236.51, 236.49, 236.46, 236.44, 236.41, 236.39, 236.36, 
    236.33, 236.3, 236.27, 236.24, 236.21, 236.18, 236.15, 236.13, 236.1, 
    236.07, 236.04, 236.01, 235.98, 235.95, 235.93, 235.9, 235.87, 235.85, 
    235.82, 235.79, 235.77, 235.74, 235.72, 235.69, 235.67, 235.64, 235.61, 
    235.58, 235.55, 235.52, 235.5, 235.47, 235.44, 235.42, 235.39, 235.36, 
    235.34, 235.31, 235.28, 235.26, 235.24, 235.21, 235.19, 235.17, 235.14, 
    235.12, 235.1, 235.07, 235.05, 235.03, 235.01, 234.98, 234.96, 234.93, 
    234.91, 234.88, 234.86, 234.84, 234.81, 234.79, 234.77, 234.74, 234.72, 
    234.7, 234.68, 234.66, 234.64, 234.62, 234.6, 234.58, 234.56, 234.54, 
    234.52, 234.5, 234.48, 234.47, 234.45, 234.43, 234.41, 234.39, 234.38, 
    234.36, 234.34, 234.32, 234.31, 234.29, 234.27, 234.26, 234.24, 234.22, 
    234.21, 234.19, 234.18, 234.16, 234.14, 234.12, 234.1, 234.09, 234.07, 
    234.05, 234.04, 234.02, 234, 233.99, 233.97, 233.95, 233.94, 233.92, 
    233.9, 233.88, 233.86, 233.84, 233.82, 233.8, 233.78, 233.75, 233.73, 
    233.71, 233.68, 233.66, 233.63, 233.6, 233.58, 233.55, 233.53, 233.5, 
    233.47, 233.44, 233.41, 233.38, 233.35, 233.33, 233.3, 233.27, 233.24, 
    233.21, 233.17, 233.14, 233.11, 233.07, 233.04, 233, 232.97, 232.93, 
    232.89, 232.85, 232.81, 232.77, 232.74, 232.7, 232.66, 232.62, 232.59, 
    232.55, 232.51, 232.47, 232.44, 232.4, 232.36, 232.33, 232.29, 232.25, 
    232.22, 232.18, 232.15, 232.11, 232.07, 232.04, 232, 231.97, 231.93, 
    231.9, 231.86, 231.83, 231.79, 231.76, 231.72, 231.69, 231.66, 231.63, 
    231.6, 231.57, 231.54, 231.51, 231.48, 231.45, 231.42, 231.39, 231.36, 
    231.34, 231.31, 231.28, 231.25, 231.22, 231.19, 231.17, 231.14, 231.11, 
    231.08, 231.05, 231.03, 231, 230.97, 230.94, 230.92, 230.89, 230.86, 
    230.84, 230.81, 230.79, 230.76, 230.74, 230.72, 230.69, 230.67, 230.65, 
    230.62, 230.6, 230.58, 230.56, 230.53, 230.51, 230.49, 230.46, 230.44, 
    230.41, 230.39, 230.37, 230.35, 230.33, 230.3, 230.28, 230.26, 230.24, 
    230.22, 230.21, 230.19, 230.17, 230.15, 230.13, 230.11, 230.09, 230.07, 
    230.05, 230.03, 230.01, 229.99, 229.97, 229.94, 229.92, 229.9, 229.88, 
    229.86, 229.84, 229.82, 229.8, 229.78, 229.76, 229.74, 229.72, 229.7, 
    229.69, 229.67, 229.65, 229.63, 229.61, 229.59, 229.58, 229.56, 229.54, 
    229.52, 229.49, 229.47, 229.45, 229.43, 229.4, 229.38, 229.36, 229.33, 
    229.31, 229.29, 229.27, 229.25, 229.23, 229.2, 229.18, 229.16, 229.14, 
    229.12, 229.1, 229.08, 229.06, 229.03, 229.01, 228.99, 228.97, 228.94, 
    228.92, 228.9, 228.88, 228.85, 228.83, 228.8, 228.78, 228.75, 228.73, 
    228.71, 228.68, 228.66, 228.64, 228.61, 228.59, 228.57, 228.55, 228.53, 
    228.51, 228.49, 228.47, 228.45, 228.43, 228.41, 228.39, 228.37, 228.35, 
    228.33, 228.31, 228.29, 228.27, 228.25, 228.23, 228.21, 228.19, 228.16, 
    228.14, 228.12, 228.1, 228.08, 228.05, 228.03, 228.01, 227.99, 227.97, 
    227.95, 227.93, 227.91, 227.89, 227.87, 227.85, 227.83, 227.81, 227.79, 
    227.77, 227.74, 227.72, 227.7, 227.67, 227.65, 227.63, 227.6, 227.58, 
    227.55, 227.53, 227.5, 227.48, 227.45, 227.43, 227.4, 227.38, 227.35, 
    227.33, 227.3, 227.28, 227.26, 227.23, 227.21, 227.19, 227.16, 227.14, 
    227.11, 227.09, 227.06, 227.03, 227.01, 226.98, 226.95, 226.93, 226.9, 
    226.88, 226.85, 226.83, 226.81, 226.78, 226.76, 226.73, 226.71, 226.68, 
    226.66, 226.64, 226.61, 226.58, 226.56, 226.53, 226.51, 226.48, 226.45, 
    226.43, 226.4, 226.38, 226.35, 226.32, 226.29, 226.27, 226.24, 226.21, 
    226.19, 226.16, 226.14, 226.11, 226.09, 226.07, 226.05, 226.02, 226, 
    225.98, 225.96, 225.94, 225.92, 225.9, 225.88, 225.85, 225.83, 225.81, 
    225.79, 225.76, 225.74, 225.72, 225.69, 225.67, 225.65, 225.63, 225.61, 
    225.58, 225.56, 225.54, 225.52, 225.49, 225.47, 225.45, 225.43, 225.41, 
    225.39, 225.37, 225.34, 225.32, 225.3, 225.28, 225.26, 225.24, 225.22, 
    225.2, 225.18, 225.15, 225.13, 225.11, 225.08, 225.05, 225.03, 225, 
    224.98, 224.95, 224.93, 224.91, 224.88, 224.86, 224.83, 224.81, 224.78, 
    224.75, 224.73, 224.7, 224.68, 224.66, 224.63, 224.61, 224.58, 224.56, 
    224.53, 224.51, 224.49, 224.46, 224.44, 224.41, 224.39, 224.36, 224.33, 
    224.31, 224.28, 224.25, 224.22, 224.19, 224.16, 224.13, 224.11, 224.08, 
    224.05, 224.02, 224, 223.97, 223.94, 223.92, 223.89, 223.86, 223.84, 
    223.81, 223.79, 223.76, 223.73, 223.7, 223.68, 223.65, 223.62, 223.59, 
    223.56, 223.53, 223.5, 223.46, 223.43, 223.4, 223.37, 223.34, 223.31, 
    223.28, 223.25, 223.22, 223.19, 223.16, 223.13, 223.1, 223.07, 223.04, 
    223.01, 222.98, 222.95, 222.92, 222.89, 222.86, 222.84, 222.81, 222.78, 
    222.75, 222.72, 222.69, 222.66, 222.63, 222.6, 222.58, 222.55, 222.53, 
    222.51, 222.48, 222.46, 222.43, 222.41, 222.39, 222.37, 222.35, 222.33, 
    222.3, 222.28, 222.25, 222.23, 222.2, 222.18, 222.15, 222.13, 222.1, 
    222.07, 222.04, 222.02, 221.99, 221.97, 221.94, 221.92, 221.89, 221.86, 
    221.83, 221.8, 221.78, 221.75, 221.72, 221.69, 221.66, 221.64, 221.61, 
    221.58, 221.55, 221.52, 221.49, 221.45, 221.42, 221.39, 221.36, 221.33, 
    221.29, 221.26, 221.23, 221.19, 221.16, 221.13, 221.09, 221.06, 221.03, 
    220.99, 220.96, 220.93, 220.9, 220.88, 220.85, 220.82, 220.79, 220.76, 
    220.73, 220.7, 220.68, 220.65, 220.62, 220.6, 220.57, 220.54, 220.52, 
    220.49, 220.46, 220.44, 220.41, 220.39, 220.36, 220.33, 220.31, 220.28, 
    220.26, 220.23, 220.21, 220.19, 220.16, 220.14, 220.12, 220.1, 220.07, 
    220.05, 220.03, 220.01, 219.99, 219.97, 219.95, 219.92, 219.9, 219.88, 
    219.86, 219.84, 219.82, 219.8, 219.78, 219.75, 219.73, 219.71, 219.69, 
    219.67, 219.64, 219.62, 219.6, 219.57, 219.55, 219.52, 219.49, 219.47, 
    219.44, 219.42, 219.39, 219.37, 219.34, 219.32, 219.29, 219.27, 219.24, 
    219.22, 219.19, 219.17, 219.14, 219.11, 219.09, 219.06, 219.04, 219.01, 
    218.99, 218.96, 218.94, 218.91, 218.88, 218.85, 218.82, 218.8, 218.77, 
    218.74, 218.71, 218.68, 218.65, 218.63, 218.6, 218.57, 218.55, 218.52, 
    218.5, 218.47, 218.44, 218.42, 218.39, 218.36, 218.34, 218.31, 218.27, 
    218.24, 218.21, 218.19, 218.16, 218.13, 218.1, 218.07, 218.05, 218.02, 
    217.99, 217.96, 217.93, 217.9, 217.87, 217.85, 217.82, 217.79, 217.76, 
    217.74, 217.71, 217.69, 217.66, 217.64, 217.62, 217.6, 217.57, 217.55, 
    217.53, 217.51, 217.49, 217.47, 217.44, 217.42, 217.4, 217.37, 217.35, 
    217.33, 217.31, 217.29, 217.27, 217.25, 217.23, 217.21, 217.19, 217.17, 
    217.15, 217.13, 217.12, 217.1, 217.08, 217.06, 217.05, 217.03, 217.01, 
    217, 216.98, 216.96, 216.94, 216.92, 216.9, 216.88, 216.86, 216.84, 
    216.81, 216.79, 216.77, 216.75, 216.72, 216.7, 216.68, 216.66, 216.64, 
    216.63, 216.61, 216.59, 216.57, 216.55, 216.53, 216.52, 216.5, 216.47, 
    216.45, 216.43, 216.41, 216.38, 216.36, 216.33, 216.3, 216.28, 216.25, 
    216.22, 216.19, 216.16, 216.13, 216.1, 216.07, 216.05, 216.02, 215.99, 
    215.96, 215.93, 215.91, 215.88, 215.85, 215.82, 215.8, 215.77, 215.74, 
    215.71, 215.68, 215.64, 215.61, 215.58, 215.54, 215.51, 215.48, 215.45, 
    215.42, 215.38, 215.35, 215.32, 215.29, 215.26, 215.23, 215.21, 215.18, 
    215.15, 215.12, 215.09, 215.06, 215.03, 215, 214.97, 214.94, 214.9, 
    214.87, 214.84, 214.81, 214.77, 214.74, 214.71, 214.67, 214.64, 214.61, 
    214.58, 214.55, 214.51, 214.48, 214.45, 214.42, 214.39, 214.36, 214.32, 
    214.29, 214.26, 214.23, 214.2, 214.16, 214.13, 214.1, 214.07, 214.04, 
    214.01, 213.98, 213.95, 213.92, 213.89, 213.86, 213.82, 213.79, 213.76, 
    213.74, 213.71, 213.68, 213.65, 213.62, 213.59, 213.57, 213.54, 213.51, 
    213.48, 213.46, 213.43, 213.4, 213.37, 213.34, 213.32, 213.29, 213.26, 
    213.24, 213.21, 213.19, 213.16, 213.13, 213.11, 213.08, 213.06, 213.03, 
    213, 212.98, 212.95, 212.92, 212.89, 212.87, 212.84, 212.81, 212.79, 
    212.77, 212.74, 212.72, 212.7, 212.67, 212.65, 212.63, 212.61, 212.58, 
    212.56, 212.54, 212.51, 212.49, 212.47, 212.45, 212.43, 212.41, 212.39, 
    212.37, 212.35, 212.33, 212.31, 212.28, 212.26, 212.24, 212.22, 212.2, 
    212.17, 212.15, 212.13, 212.1, 212.08, 212.06, 212.03, 212.01, 211.98, 
    211.96, 211.94, 211.91, 211.89, 211.86, 211.84, 211.81, 211.79, 211.76, 
    211.74, 211.71, 211.69, 211.66, 211.64, 211.61, 211.59, 211.56, 211.54, 
    211.51, 211.49, 211.46, 211.44, 211.42, 211.39, 211.37, 211.34, 211.32, 
    211.3, 211.28, 211.25, 211.23, 211.21, 211.19, 211.17, 211.15, 211.12, 
    211.1, 211.08, 211.06, 211.04, 211.02, 211, 210.97, 210.95, 210.93, 
    210.91, 210.89, 210.86, 210.84, 210.82, 210.8, 210.78, 210.75, 210.73, 
    210.71, 210.69, 210.67, 210.65, 210.63, 210.61, 210.59, 210.57, 210.54, 
    210.52, 210.5, 210.48, 210.46, 210.44, 210.42, 210.4, 210.38, 210.36, 
    210.34, 210.32, 210.3, 210.28, 210.26, 210.24, 210.22, 210.21, 210.19, 
    210.17, 210.15, 210.13, 210.12, 210.1, 210.08, 210.06, 210.04, 210.02, 
    209.99, 209.97, 209.95, 209.92, 209.9, 209.87, 209.85, 209.82, 209.8, 
    209.77, 209.75, 209.72, 209.7, 209.68, 209.66, 209.63, 209.61, 209.59, 
    209.57, 209.54, 209.52, 209.5, 209.47, 209.45, 209.43, 209.4, 209.38, 
    209.35, 209.32, 209.3, 209.27, 209.24, 209.22, 209.19, 209.16, 209.13, 
    209.11, 209.08, 209.05, 209.03, 209, 208.98, 208.96, 208.93, 208.91, 
    208.88, 208.86, 208.84, 208.81, 208.78, 208.76, 208.73, 208.7, 208.67, 
    208.64, 208.62, 208.59, 208.56, 208.54, 208.51, 208.48, 208.45, 208.43, 
    208.4, 208.38, 208.35, 208.32, 208.3, 208.27, 208.24, 208.21, 208.18, 
    208.15, 208.13, 208.1, 208.08, 208.05, 208.03, 208, 207.98, 207.95, 
    207.93, 207.91, 207.88, 207.86, 207.84, 207.81, 207.79, 207.76, 207.74, 
    207.71, 207.69, 207.66, 207.64, 207.61, 207.59, 207.56, 207.53, 207.51, 
    207.48, 207.45, 207.43, 207.4, 207.38, 207.35, 207.33, 207.31, 207.29, 
    207.27, 207.25, 207.23, 207.21, 207.19, 207.17, 207.14, 207.12, 207.1, 
    207.07, 207.05, 207.02, 207, 206.97, 206.95, 206.92, 206.9, 206.87, 
    206.85, 206.82, 206.8, 206.77, 206.74, 206.72, 206.69, 206.67, 206.65, 
    206.62, 206.6, 206.57, 206.55, 206.52, 206.5, 206.47, 206.45, 206.42, 
    206.4, 206.37, 206.34, 206.32, 206.29, 206.26, 206.24, 206.21, 206.18, 
    206.15, 206.13, 206.1, 206.08, 206.05, 206.03, 206.01, 205.98, 205.96, 
    205.93, 205.91, 205.89, 205.87, 205.85, 205.83, 205.8, 205.78, 205.76, 
    205.73, 205.71, 205.68, 205.66, 205.64, 205.62, 205.59, 205.57, 205.55, 
    205.52, 205.5, 205.48, 205.45, 205.43, 205.4, 205.38, 205.35, 205.32, 
    205.3, 205.27, 205.24, 205.21, 205.19, 205.16, 205.13, 205.1, 205.07, 
    205.04, 205.01, 204.98, 204.95, 204.92, 204.89, 204.86, 204.83, 204.8, 
    204.77, 204.74, 204.71, 204.68, 204.65, 204.61, 204.58, 204.55, 204.52, 
    204.49, 204.46, 204.42, 204.4, 204.37, 204.34, 204.31, 204.29, 204.27, 
    204.24, 204.22, 204.19, 204.17, 204.15, 204.12, 204.1, 204.07, 204.05, 
    204.03, 204.01, 203.98, 203.96, 203.94, 203.91, 203.89, 203.87, 203.85, 
    203.83, 203.81, 203.79, 203.78, 203.76, 203.74, 203.73, 203.71, 203.7, 
    203.68, 203.67, 203.66, 203.64, 203.63, 203.62, 203.6, 203.59, 203.57, 
    203.56, 203.55, 203.53, 203.52, 203.51, 203.5, 203.49, 203.48, 203.47, 
    203.46, 203.44, 203.43, 203.42, 203.41, 203.41, 203.4, 203.39, 203.39, 
    203.38, 203.37, 203.37, 203.37, 203.36, 203.36, 203.35, 203.35, 203.35, 
    203.34, 203.34, 203.33, 203.32, 203.31, 203.31, 203.3, 203.29, 203.29, 
    203.29, 203.28, 203.28, 203.27, 203.27, 203.27, 203.26, 203.26, 203.26, 
    203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 
    203.26, 203.26, 203.25, 203.25, 203.24, 203.24, 203.23, 203.23, 203.23, 
    203.22, 203.22, 203.22, 203.23, 203.23, 203.23, 203.24, 203.24, 203.24, 
    203.25, 203.25, 203.25, 203.26, 203.26, 203.27, 203.27, 203.27, 203.28, 
    203.28, 203.29, 203.3, 203.3, 203.31, 203.32, 203.32, 203.33, 203.34, 
    203.35, 203.36, 203.37, 203.38, 203.39, 203.4, 203.41, 203.43, 203.44, 
    203.45, 203.46, 203.47, 203.48, 203.5, 203.51, 203.52, 203.54, 203.55, 
    203.56, 203.58, 203.59, 203.61, 203.62, 203.64, 203.65, 203.66, 203.68, 
    203.69, 203.7, 203.71, 203.72, 203.73, 203.75, 203.76, 203.78, 203.79, 
    203.81, 203.83, 203.84, 203.86, 203.88, 203.9, 203.93, 203.95, 203.97, 
    204, 204.02, 204.04, 204.06, 204.09, 204.11, 204.13, 204.15, 204.17, 
    204.19, 204.21, 204.23, 204.24, 204.25, 204.26, 204.28, 204.29, 204.3, 
    204.31, 204.32, 204.33, 204.34, 204.34, 204.35, 204.36, 204.36, 204.36, 
    204.36, 204.35, 204.35, 204.34, 204.33, 204.32, 204.31, 204.3, 204.29, 
    204.27, 204.26, 204.24, 204.23, 204.21, 204.19, 204.17, 204.15, 204.13, 
    204.11, 204.08, 204.06, 204.04, 204.02, 204, 203.98, 203.96, 203.94, 
    203.92, 203.9, 203.88, 203.86, 203.84, 203.83, 203.81, 203.79, 203.78, 
    203.76, 203.75, 203.74, 203.73, 203.71, 203.7, 203.69, 203.67, 203.66, 
    203.65, 203.63, 203.61, 203.6, 203.58, 203.56, 203.54, 203.52, 203.5, 
    203.48, 203.47, 203.45, 203.43, 203.41, 203.39, 203.37, 203.35, 203.34, 
    203.32, 203.3, 203.28, 203.26, 203.24, 203.22, 203.2, 203.18, 203.17, 
    203.14, 203.12, 203.1, 203.08, 203.06, 203.03, 203.01, 202.99, 202.97, 
    202.95, 202.93, 202.91, 202.89, 202.88, 202.86, 202.85, 202.83, 202.82, 
    202.81, 202.79, 202.78, 202.78, 202.77, 202.76, 202.76, 202.75, 202.75, 
    202.75, 202.75, 202.75, 202.76, 202.76, 202.77, 202.78, 202.79, 202.8, 
    202.81, 202.81, 202.82, 202.83, 202.84, 202.85, 202.86, 202.87, 202.87, 
    202.88, 202.89, 202.9, 202.91, 202.92, 202.93, 202.94, 202.95, 202.96, 
    202.97, 202.98, 202.99, 203, 203.01, 203.02, 203.03, 203.04, 203.04, 
    203.05, 203.06, 203.06, 203.07, 203.07, 203.08, 203.08, 203.08, 203.09, 
    203.09, 203.09, 203.1, 203.1, 203.11, 203.11, 203.12, 203.12, 203.13, 
    203.14, 203.15, 203.16, 203.17, 203.19, 203.2, 203.22, 203.24, 203.26, 
    203.28, 203.3, 203.32, 203.34, 203.36, 203.38, 203.39, 203.41, 203.43, 
    203.45, 203.46, 203.47, 203.49, 203.5, 203.51, 203.51, 203.52, 203.53, 
    203.55, 203.56, 203.57, 203.58, 203.59, 203.6, 203.61, 203.62, 203.63, 
    203.63, 203.64, 203.65, 203.65, 203.66, 203.66, 203.66, 203.65, 203.65, 
    203.64, 203.64, 203.63, 203.63, 203.63, 203.63, 203.63, 203.63, 203.64, 
    203.64, 203.65, 203.66, 203.67, 203.69, 203.7, 203.72, 203.73, 203.75, 
    203.77, 203.79, 203.8, 203.82, 203.83, 203.85, 203.87, 203.89, 203.91, 
    203.92, 203.94, 203.96, 203.98, 204, 204.03, 204.05, 204.07, 204.09, 
    204.12, 204.14, 204.16, 204.18, 204.2, 204.21, 204.23, 204.25, 204.26, 
    204.27, 204.29, 204.3, 204.31, 204.33, 204.34, 204.36, 204.37, 204.39, 
    204.4, 204.42, 204.43, 204.45, 204.46, 204.48, 204.49, 204.51, 204.53, 
    204.54, 204.56, 204.57, 204.59, 204.61, 204.63, 204.65, 204.67, 204.69, 
    204.71, 204.73, 204.75, 204.78, 204.8, 204.83, 204.86, 204.88, 204.91, 
    204.94, 204.96, 204.99, 205.01, 205.03, 205.05, 205.07, 205.08, 205.09, 
    205.11, 205.12, 205.13, 205.14, 205.15, 205.17, 205.18, 205.19, 205.21, 
    205.22, 205.23, 205.25, 205.26, 205.28, 205.29, 205.31, 205.32, 205.33, 
    205.35, 205.36, 205.38, 205.39, 205.4, 205.42, 205.43, 205.45, 205.46, 
    205.47, 205.49, 205.5, 205.51, 205.52, 205.53, 205.54, 205.55, 205.56, 
    205.57, 205.58, 205.59, 205.6, 205.61, 205.62, 205.63, 205.63, 205.64, 
    205.64, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 
    205.65, 205.65, 205.64, 205.64, 205.63, 205.62, 205.61, 205.6, 205.58, 
    205.57, 205.56, 205.55, 205.54, 205.53, 205.51, 205.5, 205.49, 205.49, 
    205.48, 205.48, 205.48, 205.48, 205.47, 205.47, 205.48, 205.48, 205.48, 
    205.49, 205.5, 205.51, 205.52, 205.53, 205.54, 205.55, 205.55, 205.56, 
    205.57, 205.58, 205.59, 205.59, 205.6, 205.61, 205.62, 205.63, 205.64, 
    205.65, 205.66, 205.68, 205.69, 205.7, 205.72, 205.73, 205.75, 205.77, 
    205.78, 205.8, 205.81, 205.82, 205.84, 205.85, 205.87, 205.88, 205.89, 
    205.91, 205.92, 205.93, 205.94, 205.94, 205.95, 205.96, 205.97, 205.98, 
    205.99, 206, 206.01, 206.02, 206.04, 206.05, 206.07, 206.08, 206.1, 
    206.12, 206.13, 206.15, 206.17, 206.19, 206.21, 206.23, 206.25, 206.26, 
    206.28, 206.3, 206.31, 206.33, 206.34, 206.36, 206.37, 206.39, 206.4, 
    206.41, 206.43, 206.44, 206.45, 206.46, 206.47, 206.48, 206.49, 206.49, 
    206.5, 206.5, 206.5, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 
    206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 
    206.51, 206.51, 206.52, 206.52, 206.52, 206.52, 206.52, 206.52, 206.53, 
    206.53, 206.53, 206.53, 206.53, 206.53, 206.54, 206.54, 206.54, 206.54, 
    206.55, 206.55, 206.56, 206.57, 206.58, 206.59, 206.6, 206.61, 206.62, 
    206.63, 206.64, 206.66, 206.67, 206.68, 206.69, 206.7, 206.71, 206.71, 
    206.72, 206.73, 206.73, 206.74, 206.75, 206.76, 206.77, 206.78, 206.79, 
    206.8, 206.81, 206.83, 206.84, 206.85, 206.87, 206.88, 206.89, 206.9, 
    206.91, 206.92, 206.93, 206.94, 206.95, 206.96, 206.97, 206.98, 206.99, 
    207, 207, 207.01, 207.02, 207.03, 207.03, 207.04, 207.04, 207.05, 207.05, 
    207.06, 207.06, 207.07, 207.07, 207.07, 207.07, 207.08, 207.08, 207.07, 
    207.07, 207.07, 207.06, 207.06, 207.06, 207.05, 207.05, 207.04, 207.04, 
    207.03, 207.03, 207.03, 207.02, 207.02, 207.02, 207.02, 207.02, 207.02, 
    207.02, 207.01, 207.01, 207, 207, 206.99, 206.98, 206.97, 206.95, 206.96, 
    206.97, 206.98, 206.99, 207, 207.01, 207.02, 207.03, 207.04, 207.04, 
    207.05, 207.05, 207.06, 207.06, 207.06, 207.06, 207.06, 207.05, 207.05, 
    207.04, 207.03, 207.02, 207.01, 207, 206.99, 206.97, 206.96, 206.95, 
    206.94, 206.92, 206.91, 206.9, 206.9, 206.89, 206.88, 206.88, 206.87, 
    206.87, 206.87, 206.86, 206.86, 206.86, 206.86, 206.86, 206.86, 206.86, 
    206.86, 206.86, 206.86, 206.85, 206.85, 206.85, 206.85, 206.84, 206.84, 
    206.84, 206.83, 206.83, 206.82, 206.82, 206.81, 206.81, 206.81, 206.8, 
    206.8, 206.8, 206.79, 206.79, 206.79, 206.79, 206.79, 206.79, 206.8, 
    206.8, 206.8, 206.8, 206.81, 206.81, 206.81, 206.82, 206.82, 206.82, 
    206.82, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 
    206.83, 206.83, 206.83, 206.82, 206.82, 206.82, 206.82, 206.81, 206.81, 
    206.81, 206.8, 206.8, 206.8, 206.8, 206.79, 206.79, 206.79, 206.78, 
    206.78, 206.78, 206.78, 206.77, 206.77, 206.77, 206.77, 206.77, 206.76, 
    206.76, 206.76, 206.76, 206.76, 206.75, 206.75, 206.75, 206.75, 206.74, 
    206.74, 206.74, 206.73, 206.73, 206.73, 206.72, 206.72, 206.71, 206.7, 
    206.69, 206.69, 206.68, 206.67, 206.65, 206.64, 206.63, 206.61, 206.6, 
    206.58, 206.56, 206.54, 206.52, 206.49, 206.47, 206.44, 206.41, 206.39, 
    206.36, 206.32, 206.29, 206.26, 206.23, 206.19, 206.16, 206.12, 206.09, 
    206.05, 206.02, 205.98, 205.94, 205.91, 205.87, 205.83, 205.8, 205.76, 
    205.73, 205.69, 205.65, 205.62, 205.58, 205.55, 205.51, 205.48, 205.44, 
    205.41, 205.37, 205.33, 205.3, 205.26, 205.23, 205.19, 205.16, 205.12, 
    205.08, 205.05, 205.01, 204.97, 204.93, 204.89, 204.86, 204.82, 204.77, 
    204.73, 204.69, 204.65, 204.6, 204.55, 204.5, 204.45, 204.4, 204.35, 
    204.29, 204.23, 204.17, 204.11, 204.05, 203.98, 203.91, 203.84, 203.77, 
    203.7, 203.62, 203.55, 203.47, 203.4, 203.32, 203.25, 203.17, 203.1, 
    203.03, 202.96, 202.89, 202.82, 202.75, 202.69, 202.63, 202.57, 202.51, 
    202.45, 202.4, 202.35, 202.3, 202.25, 202.21, 202.16, 202.12, 202.08, 
    202.05, 202.01, 201.98, 201.95, 201.93, 201.9, 201.88, 201.87, 201.85, 
    201.84, 201.83, 201.82, 201.82, 201.82, 201.82, 201.82, 201.83, 201.84, 
    201.85, 201.86, 201.87, 201.88, 201.9, 201.91, 201.93, 201.95, 201.96, 
    201.98, 201.99, 202.01, 202.02, 202.04, 202.05, 202.06, 202.07, 202.08, 
    202.09, 202.09, 202.1, 202.1, 202.1, 202.1, 202.1, 202.1, 202.1, 202.09, 
    202.09, 202.08, 202.07, 202.06, 202.05, 202.04, 202.03, 202.01, 201.99, 
    201.97, 201.95, 201.93, 201.9, 201.87, 201.84, 201.81, 201.77, 201.73, 
    201.69, 201.65, 201.6, 201.55, 201.5, 201.44, 201.39, 201.33, 201.27, 
    201.2, 201.14, 201.07, 201.01, 200.94, 200.87, 200.8, 200.73, 200.65, 
    200.58, 200.51, 200.44, 200.37, 200.29, 200.22, 200.15, 200.09, 200.02, 
    199.95, 199.89, 199.83, 199.77, 199.71, 199.65, 199.6, 199.55, 199.5, 
    199.46, 199.42, 199.38, 199.34, 199.31, 199.28, 199.25, 199.23, 199.21, 
    199.19, 199.18, 199.16, 199.15, 199.15, 199.14, 199.14, 199.14, 199.15, 
    199.15, 199.16, 199.17, 199.18, 199.19, 199.21, 199.22, 199.24, 199.26, 
    199.28, 199.3, 199.32, 199.35, 199.37, 199.39, 199.42, 199.44, 199.47, 
    199.49, 199.52, 199.55, 199.57, 199.6, 199.62, 199.65, 199.67, 199.7, 
    199.72, 199.75, 199.77, 199.8, 199.82, 199.84, 199.86, 199.88, 199.9, 
    199.91, 199.93, 199.94, 199.95, 199.96, 199.97, 199.98, 199.98, 199.98, 
    199.98, 199.98, 199.98, 199.97, 199.97, 199.96, 199.96, 199.95, 199.94, 
    199.93, 199.93, 199.92, 199.91, 199.91, 199.91, 199.9, 199.9, 199.9, 
    199.9, 199.9, 199.91, 199.91, 199.92, 199.92, 199.93, 199.94, 199.95, 
    199.96, 199.97, 199.98, 199.98, 199.99, 200, 200.01, 200.01, 200.02, 
    200.03, 200.03, 200.03, 200.04, 200.04, 200.04, 200.04, 200.04, 200.04, 
    200.04, 200.04, 200.04, 200.03, 200.03, 200.02, 200.01, 200, 199.99, 
    199.98, 199.96, 199.95, 199.93, 199.91, 199.88, 199.86, 199.83, 199.81, 
    199.78, 199.75, 199.72, 199.69, 199.66, 199.63, 199.6, 199.57, 199.54, 
    199.52, 199.49, 199.47, 199.46, 199.44, 199.43, 199.43, 199.42, 199.42, 
    199.43, 199.44, 199.45, 199.47, 199.49, 199.52, 199.54, 199.58, 199.61, 
    199.65, 199.69, 199.73, 199.78, 199.82, 199.87, 199.92, 199.96, 200.01, 
    200.06, 200.1, 200.14, 200.18, 200.22, 200.26, 200.29, 200.31, 200.33, 
    200.35, 200.36, 200.37, 200.37, 200.37, 200.36, 200.35, 200.33, 200.31, 
    200.28, 200.25, 200.21, 200.17, 200.13, 200.09, 200.04, 199.99, 199.94, 
    199.89, 199.84, 199.8, 199.75, 199.7, 199.66, 199.62, 199.58, 199.54, 
    199.51, 199.48, 199.45, 199.43, 199.4, 199.39, 199.37, 199.36, 199.35, 
    199.34, 199.34, 199.34, 199.34, 199.35, 199.35, 199.36, 199.38, 199.4, 
    199.42, 199.44, 199.47, 199.5, 199.54, 199.58, 199.62, 199.67, 199.72, 
    199.78, 199.84, 199.91, 199.97, 200.04, 200.12, 200.19, 200.26, 200.34, 
    200.42, 200.49, 200.57, 200.64, 200.72, 200.79, 200.85, 200.92, 200.98, 
    201.04, 201.09, 201.14, 201.18, 201.22, 201.26, 201.29, 201.31, 201.33, 
    201.35, 201.36, 201.37, 201.37, 201.36, 201.36, 201.34, 201.33, 201.3, 
    201.28, 201.25, 201.22, 201.19, 201.15, 201.11, 201.07, 201.03, 200.99, 
    200.95, 200.91, 200.88, 200.84, 200.81, 200.78, 200.75, 200.73, 200.7, 
    200.69, 200.67, 200.66, 200.66, 200.65, 200.66, 200.66, 200.67, 200.68, 
    200.69, 200.71, 200.73, 200.76, 200.79, 200.82, 200.86, 200.9, 200.94, 
    200.99, 201.04, 201.09, 201.15, 201.21, 201.27, 201.33, 201.39, 201.46, 
    201.53, 201.6, 201.67, 201.75, 201.83, 201.9, 201.98, 202.07, 202.15, 
    202.24, 202.33, 202.42, 202.52, 202.61, 202.71, 202.82, 202.92, 203.02, 
    203.13, 203.23, 203.34, 203.44, 203.54, 203.64, 203.73, 203.82, 203.9, 
    203.98, 204.05, 204.11, 204.17, 204.22, 204.26, 204.29, 204.31, 204.33, 
    204.33, 204.33, 204.32, 204.3, 204.27, 204.24, 204.2, 204.15, 204.09, 
    204.03, 203.97, 203.9, 203.83, 203.75, 203.68, 203.6, 203.53, 203.45, 
    203.38, 203.32, 203.26, 203.2, 203.15, 203.11, 203.08, 203.06, 203.04, 
    203.03, 203.04, 203.05, 203.07, 203.1, 203.14, 203.18, 203.24, 203.3, 
    203.37, 203.45, 203.53, 203.62, 203.71, 203.81, 203.92, 204.03, 204.14, 
    204.26, 204.38, 204.5, 204.63, 204.76, 204.89, 205.02, 205.16, 205.29, 
    205.43, 205.57, 205.71, 205.86, 206, 206.15, 206.29, 206.44, 206.59, 
    206.74, 206.9, 207.05, 207.21, 207.36, 207.52, 207.68, 207.85, 208.01, 
    208.18, 208.35, 208.52, 208.69, 208.87, 209.05, 209.23, 209.41, 209.59, 
    209.77, 209.96, 210.15, 210.33, 210.52, 210.71, 210.9, 211.08, 211.26, 
    211.44, 211.62, 211.8, 211.96, 212.13, 212.29, 212.44, 212.58, 212.72, 
    212.84, 212.96, 213.08, 213.18, 213.28, 213.36, 213.44, 213.51, 213.58, 
    213.64, 213.69, 213.74, 213.79, 213.84, 213.88, 213.92, 213.96, 214.01, 
    214.05, 214.1, 214.15, 214.21, 214.27, 214.33, 214.4, 214.47, 214.55, 
    214.63, 214.72, 214.81, 214.91, 215.01, 215.11, 215.22, 215.33, 215.45, 
    215.56, 215.68, 215.79, 215.91, 216.03, 216.14, 216.26, 216.37, 216.48, 
    216.59, 216.69, 216.79, 216.88, 216.98, 217.06, 217.14, 217.22, 217.3, 
    217.36, 217.43, 217.49, 217.55, 217.61, 217.66, 217.72, 217.77, 217.82, 
    217.88, 217.93, 217.98, 218.04, 218.1, 218.16, 218.22, 218.28, 218.34, 
    218.41, 218.47, 218.54, 218.61, 218.68, 218.74, 218.81, 218.88, 218.94, 
    219.01, 219.07, 219.14, 219.2, 219.26, 219.33, 219.39, 219.45, 219.52, 
    219.58, 219.65, 219.72, 219.79, 219.87, 219.95, 220.04, 220.13, 220.23, 
    220.33, 220.44, 220.55, 220.67, 220.8, 220.94, 221.09, 221.24, 221.4, 
    221.56, 221.74, 221.92, 222.1, 222.29, 222.49, 222.69, 222.89, 223.1, 
    223.31, 223.53, 223.74, 223.96, 224.18, 224.4, 224.62, 224.84, 225.06, 
    225.28, 225.5, 225.71, 225.93, 226.14, 226.35, 226.56, 226.77, 226.97, 
    227.17, 227.36, 227.55, 227.74, 227.92, 228.1, 228.27, 228.43, 228.6, 
    228.75, 228.91, 229.06, 229.2, 229.35, 229.49, 229.63, 229.77, 229.91, 
    230.05, 230.2, 230.35, 230.5, 230.65, 230.81, 230.97, 231.13, 231.3, 
    231.47, 231.64, 231.81, 231.98, 232.15, 232.32, 232.48, 232.64, 232.8, 
    232.95, 233.09, 233.23, 233.37, 233.5, 233.62, 233.74, 233.85, 233.97, 
    234.07, 234.18, 234.28, 234.39, 234.49, 234.6, 234.71, 234.82, 234.94, 
    235.06, 235.19, 235.33, 235.47, 235.62, 235.78, 235.95, 236.13, 236.32, 
    236.51, 236.72, 236.93, 237.15, 237.38, 237.61, 237.86, 238.11, 238.36, 
    238.62, 238.88, 239.15, 239.42, 239.69, 239.96, 240.24, 240.5, 240.77, 
    241.04, 241.3, 241.55, 241.8, 242.05, 242.28, 242.51, 242.73, 242.95, 
    243.15, 243.34, 243.53, 243.71, 243.87, 244.03, 244.18, 244.33, 244.46, 
    244.59, 244.71, 244.82, 244.93, 245.03, 245.13, 245.23, 245.32, 245.42, 
    245.51, 245.61, 245.71, 245.81, 245.91, 246.02, 246.13, 246.25, 246.37, 
    246.5, 246.64, 246.78, 246.93, 247.09, 247.25, 247.42, 247.6, 247.78, 
    247.96, 248.15, 248.35, 248.55, 248.75, 248.96, 249.17, 249.38, 249.6, 
    249.82, 250.04, 250.26, 250.49, 250.72, 250.95, 251.18, 251.42, 251.65, 
    251.89, 252.13, 252.36, 252.6, 252.84, 253.07, 253.31, 253.55, 253.78, 
    254.01, 254.25, 254.48, 254.71, 254.93, 255.16, 255.38, 255.61, 255.83, 
    256.05, 256.27, 256.49, 256.71, 256.92, 257.14, 257.36, 257.57, 257.79, 
    258, 258.21, 258.43, 258.64, 258.85, 259.06, 259.27, 259.48, 259.69, 
    259.9, 260.11, 260.32, 260.52, 260.73, 260.94, 261.14, 261.35, 261.56, 
    261.77, 261.98, 262.19, 262.4, 262.61, 262.83, 263.04, 263.26, 263.48, 
    263.7, 263.92, 264.14, 264.36, 264.59, 264.81, 265.04, 265.26, 265.49, 
    265.72, 265.95, 266.17, 266.4, 266.63, 266.86, 267.09, 267.32, 267.55, 
    267.77, 268, 268.22, 268.45, 268.67, 268.89, 269.11, 269.32, 269.53, 
    269.75, 269.95, 270.16, 270.36, 270.56, 270.76, 270.96, 271.15, 271.34, 
    271.53, 271.71, 271.9, 272.08, 272.26, 272.44, 272.62, 272.8, 272.98, 
    273.16, 273.33, 273.51, 273.68, 273.86, 274.04, 274.21, 274.39, 274.57, 
    274.74, 274.92, 275.1, 275.27, 275.45, 275.63, 275.81, 275.99, 276.17, 
    276.35, 276.52, 276.7, 276.88, 277.06, 277.23, 277.41, 277.58, 277.75, 
    277.92, 278.08, 278.25, 278.41, 278.57, 278.72, 278.88, 279.03, 279.18, 
    279.32, 279.47, 279.61, 279.75, 279.9, 280.04, 280.18, 280.33, 280.48, 
    280.63, 280.79, 280.95, 281.11, 281.28, 281.45, 281.63, 281.81, 281.99, 
    282.18, 282.37, 282.57, 282.76, 282.96, 283.16, 283.36, 283.55, 283.75, 
    283.94, 284.13, 284.32, 284.5, 284.68, 284.86, 285.02, 285.19, 285.35, 
    285.5, 285.65, 285.79, 285.92, 286.05, 286.18, 286.3, 286.41, 286.52, 
    286.62, 286.72, 286.82, 286.91, 287, 287.09, 287.18, 287.26, 287.35, 
    287.43, 287.51, 287.6, 287.68, 287.77, 287.86, 287.95, 288.04, 288.14, 
    288.24, 288.33, 288.44, 288.54, 288.65, 288.75, 288.86, 288.97, 289.09, 
    289.2, 289.31, 289.42, 289.53, 289.65, 289.76, 289.86, 289.97, 290.07, 
    290.17, 290.27, 290.37, 290.46, 290.55, 290.63, 290.71, 290.78, 290.85, 
    290.92, 290.98, 291.04, 291.09, 291.14, 291.18, 291.22, 291.25, 291.28, 
    291.31, 291.33, 291.34, 291.35, 291.35, 291.35, 291.34, 291.32, 291.3, 
    291.27, 291.23, 291.19, 291.14, 291.08, 291.01, 290.93, 290.83, 290.72, 
    290.59, 290.46, 290.33, 290.19, 290.05, 289.91, 289.77, 289.62, 289.48, 
    289.34, 289.19, 289.05, 288.91, 288.76, 288.62, 288.48, 288.34, 288.2, 
    288.06, 287.92, 287.79, 287.65, 287.51, 287.38, 287.24, 287.11, 286.97, 
    286.84, 286.7, 286.57, 286.43, 286.3, 286.16, 286.02, 285.89, 285.75, 
    285.62, 285.48, 285.34, 285.21, 285.07, 284.93, 284.8, 284.66, 284.53, 
    284.39, 284.26, 284.12, 283.99, 283.85, 283.72, 283.58, 283.45, 283.31, 
    283.17, 283.03, 282.9, 282.76, 282.62, 282.47, 282.33, 282.19, 282.04, 
    281.9, 281.75, 281.6, 281.45, 281.3, 281.15, 281, 280.85, 280.7, 280.55, 
    280.39, 280.24, 280.09, 279.94, 279.79, 279.63, 279.48, 279.33, 279.17, 
    279.02, 278.86, 278.71, 278.55, 278.39, 278.23, 278.07, 277.91, 277.74, 
    277.58, 277.41, 277.24, 277.08, 276.91, 276.73, 276.56, 276.39, 276.22, 
    276.04, 275.87, 275.69, 275.51, 275.33, 275.15, 274.97, 274.79, 274.61, 
    274.43, 274.24, 274.06, 273.87, 273.69, 273.5, 273.31, 273.12, 272.93, 
    272.74, 272.55, 272.35, 272.16, 271.97, 271.78, 271.59, 271.4, 271.2, 
    271.01, 270.82, 270.64, 270.45, 270.26, 270.07, 269.88, 269.7, 269.51, 
    269.32, 269.13, 268.95, 268.76, 268.57, 268.38, 268.19, 268, 267.81, 
    267.62, 267.43, 267.24, 267.05, 266.85, 266.66, 266.47, 266.27, 266.08, 
    265.88, 265.69, 265.49, 265.29, 265.1, 264.9, 264.7, 264.5, 264.31, 
    264.11, 263.91, 263.71, 263.51, 263.31, 263.11, 262.91, 262.71, 262.51, 
    262.3, 262.1, 261.9, 261.7, 261.5, 261.29, 261.09, 260.89, 260.69, 
    260.48, 260.28, 260.08, 259.87, 259.67, 259.47, 259.26, 259.06, 258.86, 
    258.65, 258.45, 258.25, 258.04, 257.84, 257.63, 257.42, 257.22, 257.01, 
    256.8, 256.59, 256.38, 256.16, 255.95, 255.74, 255.52, 255.3, 255.09, 
    254.87, 254.65, 254.43, 254.21, 253.99, 253.77, 253.55, 253.34, 253.12, 
    252.9, 252.69, 252.47, 252.26, 252.05, 251.84, 251.63, 251.43, 251.22, 
    251.02, 250.82, 250.61, 250.41, 250.22, 250.02, 249.82, 249.62, 249.43, 
    249.23, 249.04, 248.84, 248.65, 248.46, 248.26, 248.07, 247.88, 247.68, 
    247.49, 247.3, 247.11, 246.92, 246.73, 246.54, 246.35, 246.16, 245.97, 
    245.78, 245.59, 245.41, 245.22, 245.04, 244.85, 244.67, 244.49, 244.31, 
    244.13, 243.95, 243.77, 243.59, 243.41, 243.24, 243.06, 242.89, 242.72, 
    242.55, 242.38, 242.21, 242.05, 241.88, 241.72, 241.56, 241.4, 241.24, 
    241.09, 240.94, 240.79, 240.64, 240.5, 240.36, 240.23, 240.1, 239.97, 
    239.85, 239.74, 239.63 ;

 dry_temp_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 dry_temp_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 geop =
  31.017, 32.515, 33.964, 35.36, 36.725, 38.09, 39.472, 40.889, 42.331, 
    43.799, 45.325, 46.934, 48.636, 50.438, 52.35, 54.39, 56.578, 58.889, 
    61.33, 63.893, 66.584, 69.407, 72.337, 75.365, 78.42, 81.509, 84.638, 
    87.821, 91.059, 94.324, 97.614, 100.92, 104.27, 107.67, 111.12, 114.65, 
    118.24, 121.9, 125.62, 129.38, 133.19, 137.02, 140.9, 144.82, 148.76, 
    152.72, 156.67, 160.61, 164.52, 168.43, 172.33, 176.23, 180.12, 183.99, 
    187.85, 191.68, 195.5, 199.3, 203.07, 206.84, 210.64, 214.45, 218.29, 
    222.17, 226.06, 229.95, 233.82, 237.68, 241.54, 245.4, 249.26, 253.1, 
    256.93, 260.72, 264.48, 268.2, 271.91, 275.6, 279.3, 282.98, 286.65, 
    290.29, 293.9, 297.52, 301.16, 304.83, 308.51, 312.2, 315.91, 319.63, 
    323.35, 327.08, 330.84, 334.61, 338.41, 342.23, 346.05, 349.89, 353.74, 
    357.6, 361.47, 365.34, 369.22, 373.1, 376.98, 380.88, 384.79, 388.7, 
    392.63, 396.55, 400.47, 404.39, 408.32, 412.26, 416.21, 420.16, 424.1, 
    428.05, 431.99, 435.92, 439.83, 443.72, 447.6, 451.47, 455.32, 459.17, 
    463, 466.82, 470.63, 474.44, 478.25, 482.06, 485.86, 489.65, 493.45, 
    497.26, 501.06, 504.88, 508.7, 512.53, 516.36, 520.19, 524.02, 527.85, 
    531.69, 535.53, 539.36, 543.18, 547.02, 550.85, 554.69, 558.53, 562.36, 
    566.18, 570.01, 573.86, 577.72, 581.58, 585.45, 589.35, 593.27, 597.22, 
    601.21, 605.21, 609.24, 613.29, 617.37, 621.46, 625.58, 629.71, 633.88, 
    638.07, 642.29, 646.53, 650.78, 655.05, 659.34, 663.65, 667.99, 672.37, 
    676.78, 681.24, 685.73, 690.28, 694.89, 699.58, 704.36, 709.23, 714.18, 
    719.23, 724.39, 729.67, 735, 740.38, 745.76, 751.14, 756.52, 761.89, 
    767.25, 772.56, 777.83, 783.05, 788.28, 793.51, 798.75, 803.99, 809.24, 
    814.51, 819.79, 825.05, 830.3, 835.55, 840.8, 846.06, 851.3, 856.5, 
    861.61, 866.66, 871.66, 876.63, 881.56, 886.45, 891.28, 896.05, 900.72, 
    905.3, 909.77, 914.12, 918.36, 922.52, 926.61, 930.63, 934.63, 938.63, 
    942.66, 946.7, 950.76, 954.85, 958.99, 963.17, 967.38, 971.57, 975.73, 
    979.84, 983.94, 988.02, 992.07, 996.08, 1000.1, 1004, 1007.9, 1011.8, 
    1015.6, 1019.3, 1023.1, 1027, 1030.8, 1034.7, 1038.5, 1042.3, 1046.1, 
    1049.8, 1053.4, 1057.1, 1060.7, 1064.3, 1067.9, 1071.4, 1075, 1078.5, 
    1081.9, 1085.4, 1088.8, 1092.2, 1095.5, 1098.9, 1102.1, 1105.4, 1108.5, 
    1111.7, 1114.9, 1118, 1121.2, 1124.3, 1127.4, 1130.5, 1133.6, 1136.7, 
    1139.9, 1143, 1146.2, 1149.4, 1152.6, 1155.8, 1159, 1162.2, 1165.4, 
    1168.6, 1171.8, 1175, 1178.4, 1181.7, 1185.1, 1188.5, 1192, 1195.4, 
    1198.9, 1202.4, 1205.9, 1209.4, 1212.9, 1216.4, 1219.9, 1223.4, 1226.9, 
    1230.4, 1233.8, 1237.3, 1240.8, 1244.2, 1247.7, 1251.1, 1254.6, 1258.1, 
    1261.6, 1265.2, 1268.7, 1272.3, 1275.8, 1279.4, 1282.9, 1286.4, 1289.8, 
    1293.3, 1296.7, 1300.1, 1303.5, 1306.8, 1310.1, 1313.4, 1316.6, 1319.7, 
    1322.9, 1326, 1329.1, 1332.2, 1335.4, 1338.5, 1341.7, 1344.8, 1348, 
    1351.2, 1354.5, 1357.7, 1361, 1364.2, 1367.5, 1370.9, 1374.2, 1377.5, 
    1380.8, 1384.1, 1387.4, 1390.6, 1393.9, 1397.1, 1400.3, 1403.6, 1406.9, 
    1410.2, 1413.5, 1416.9, 1420.2, 1423.6, 1427.1, 1430.5, 1434, 1437.5, 
    1441, 1444.5, 1448.1, 1451.7, 1455.3, 1458.9, 1462.5, 1466.1, 1469.7, 
    1473.3, 1476.9, 1480.5, 1484.1, 1487.7, 1491.3, 1494.9, 1498.6, 1502.2, 
    1505.9, 1509.5, 1513.2, 1516.8, 1520.5, 1524.1, 1527.8, 1531.4, 1535, 
    1538.7, 1542.3, 1545.9, 1549.5, 1553, 1556.6, 1560.2, 1563.8, 1567.3, 
    1570.9, 1574.4, 1578, 1581.6, 1585.1, 1588.7, 1592.3, 1595.8, 1599.4, 
    1602.9, 1606.5, 1610, 1613.6, 1617.1, 1620.7, 1624.2, 1627.7, 1631.2, 
    1634.7, 1638.2, 1641.8, 1645.3, 1648.8, 1652.3, 1655.8, 1659.3, 1662.9, 
    1666.4, 1670, 1673.6, 1677.1, 1680.7, 1684.3, 1687.8, 1691.4, 1695, 
    1698.5, 1702.1, 1705.6, 1709.2, 1712.7, 1716.3, 1719.8, 1723.3, 1726.9, 
    1730.4, 1733.9, 1737.4, 1740.9, 1744.5, 1748, 1751.6, 1755.1, 1758.7, 
    1762.2, 1765.8, 1769.3, 1772.8, 1776.4, 1779.9, 1783.4, 1786.9, 1790.4, 
    1793.8, 1797.3, 1800.7, 1804.2, 1807.6, 1811.1, 1814.5, 1818, 1821.5, 
    1825, 1828.5, 1832, 1835.5, 1839.1, 1842.6, 1846.2, 1849.8, 1853.3, 
    1856.9, 1860.5, 1864.1, 1867.7, 1871.2, 1874.8, 1878.4, 1882, 1885.5, 
    1889.1, 1892.6, 1896.2, 1899.8, 1903.4, 1906.9, 1910.5, 1914.1, 1917.7, 
    1921.3, 1924.9, 1928.5, 1932.2, 1935.8, 1939.4, 1943.1, 1946.7, 1950.3, 
    1954, 1957.6, 1961.2, 1964.9, 1968.5, 1972.1, 1975.7, 1979.3, 1982.9, 
    1986.6, 1990.2, 1993.8, 1997.4, 2001, 2004.7, 2008.3, 2011.9, 2015.5, 
    2019.2, 2022.8, 2026.4, 2030.1, 2033.7, 2037.3, 2040.9, 2044.5, 2048.2, 
    2051.8, 2055.4, 2059, 2062.6, 2066.2, 2069.8, 2073.4, 2077, 2080.7, 
    2084.2, 2087.8, 2091.4, 2095, 2098.6, 2102.2, 2105.8, 2109.4, 2113, 
    2116.5, 2120.1, 2123.7, 2127.3, 2130.9, 2134.5, 2138.1, 2141.7, 2145.3, 
    2148.9, 2152.5, 2156.2, 2159.8, 2163.5, 2167.1, 2170.8, 2174.4, 2178.1, 
    2181.8, 2185.4, 2189.1, 2192.8, 2196.5, 2200.2, 2203.8, 2207.5, 2211.2, 
    2214.9, 2218.5, 2222.2, 2225.9, 2229.6, 2233.3, 2236.9, 2240.6, 2244.3, 
    2248, 2251.7, 2255.4, 2259.1, 2262.8, 2266.4, 2270.1, 2273.8, 2277.4, 
    2281.1, 2284.7, 2288.3, 2291.9, 2295.6, 2299.1, 2302.7, 2306.3, 2309.9, 
    2313.5, 2317, 2320.6, 2324.2, 2327.7, 2331.3, 2334.8, 2338.4, 2342, 
    2345.5, 2349.1, 2352.7, 2356.3, 2359.9, 2363.5, 2367, 2370.6, 2374.2, 
    2377.8, 2381.4, 2385, 2388.6, 2392.2, 2395.7, 2399.3, 2402.8, 2406.4, 
    2409.9, 2413.4, 2417, 2420.5, 2424.1, 2427.6, 2431.1, 2434.6, 2438.2, 
    2441.7, 2445.2, 2448.7, 2452.3, 2455.8, 2459.3, 2462.8, 2466.4, 2469.9, 
    2473.4, 2476.9, 2480.5, 2484, 2487.5, 2491, 2494.6, 2498.1, 2501.5, 2505, 
    2508.5, 2512, 2515.4, 2518.9, 2522.4, 2525.8, 2529.3, 2532.8, 2536.3, 
    2539.8, 2543.3, 2546.8, 2550.3, 2553.9, 2557.4, 2561, 2564.6, 2568.2, 
    2571.8, 2575.5, 2579.1, 2582.7, 2586.4, 2590, 2593.7, 2597.4, 2601, 
    2604.7, 2608.4, 2612.1, 2615.7, 2619.4, 2623.1, 2626.7, 2630.3, 2634, 
    2637.6, 2641.3, 2644.9, 2648.6, 2652.2, 2655.9, 2659.6, 2663.2, 2666.8, 
    2670.5, 2674.1, 2677.8, 2681.4, 2685, 2688.7, 2692.3, 2695.9, 2699.5, 
    2703.1, 2706.7, 2710.3, 2713.9, 2717.5, 2721, 2724.6, 2728.2, 2731.7, 
    2735.3, 2738.8, 2742.3, 2745.9, 2749.4, 2752.9, 2756.4, 2760, 2763.5, 
    2767, 2770.5, 2774.1, 2777.6, 2781.1, 2784.6, 2788.1, 2791.7, 2795.2, 
    2798.7, 2802.2, 2805.7, 2809.2, 2812.8, 2816.2, 2819.7, 2823.2, 2826.7, 
    2830.2, 2833.7, 2837.2, 2840.8, 2844.3, 2847.9, 2851.5, 2855.1, 2858.8, 
    2862.5, 2866.2, 2869.9, 2873.6, 2877.3, 2881.1, 2884.9, 2888.7, 2892.5, 
    2896.3, 2900.2, 2904.1, 2907.9, 2911.8, 2915.8, 2919.7, 2923.7, 2927.7, 
    2931.7, 2935.7, 2939.7, 2943.8, 2947.8, 2951.9, 2956.1, 2960.2, 2964.4, 
    2968.6, 2972.8, 2977, 2981.3, 2985.5, 2989.8, 2994.1, 2998.4, 3002.7, 
    3007, 3011.2, 3015.5, 3019.8, 3024.1, 3028.5, 3032.8, 3037.1, 3041.4, 
    3045.7, 3049.9, 3054.2, 3058.5, 3062.8, 3067.1, 3071.4, 3075.7, 3080, 
    3084.2, 3088.5, 3092.7, 3096.9, 3101.1, 3105.3, 3109.5, 3113.6, 3117.8, 
    3121.9, 3126, 3130, 3134.1, 3138.1, 3142.1, 3146, 3150, 3153.9, 3157.7, 
    3161.6, 3165.4, 3169.2, 3172.9, 3176.7, 3180.4, 3184.1, 3187.7, 3191.4, 
    3195.1, 3198.7, 3202.3, 3205.9, 3209.5, 3213.1, 3216.7, 3220.2, 3223.8, 
    3227.3, 3230.9, 3234.4, 3237.9, 3241.5, 3245, 3248.5, 3252, 3255.6, 
    3259.1, 3262.6, 3266.2, 3269.7, 3273.3, 3276.8, 3280.4, 3283.9, 3287.5, 
    3291.1, 3294.6, 3298.2, 3301.8, 3305.3, 3308.9, 3312.5, 3316, 3319.6, 
    3323.2, 3326.7, 3330.3, 3333.9, 3337.4, 3341, 3344.5, 3348, 3351.6, 
    3355.1, 3358.7, 3362.2, 3365.7, 3369.3, 3372.8, 3376.4, 3379.9, 3383.4, 
    3387, 3390.5, 3394, 3397.6, 3401.1, 3404.6, 3408.1, 3411.6, 3415.1, 
    3418.6, 3422.1, 3425.6, 3429.1, 3432.6, 3436.1, 3439.5, 3443, 3446.4, 
    3449.9, 3453.3, 3456.8, 3460.2, 3463.7, 3467.1, 3470.5, 3473.9, 3477.4, 
    3480.8, 3484.2, 3487.7, 3491.1, 3494.5, 3498, 3501.4, 3504.8, 3508.2, 
    3511.7, 3515.1, 3518.5, 3521.9, 3525.3, 3528.7, 3532.1, 3535.5, 3538.9, 
    3542.3, 3545.8, 3549.2, 3552.6, 3556, 3559.4, 3562.8, 3566.2, 3569.6, 
    3573.1, 3576.5, 3579.9, 3583.3, 3586.8, 3590.2, 3593.6, 3597, 3600.4, 
    3603.8, 3607.2, 3610.6, 3614, 3617.4, 3620.8, 3624.2, 3627.5, 3630.9, 
    3634.3, 3637.7, 3641.1, 3644.5, 3648, 3651.4, 3654.8, 3658.2, 3661.6, 
    3665, 3668.4, 3671.8, 3675.3, 3678.7, 3682.1, 3685.5, 3688.9, 3692.4, 
    3695.8, 3699.2, 3702.6, 3706.1, 3709.5, 3712.9, 3716.4, 3719.8, 3723.3, 
    3726.7, 3730.2, 3733.6, 3737.1, 3740.6, 3744.1, 3747.6, 3751, 3754.5, 
    3758, 3761.5, 3765, 3768.5, 3772, 3775.5, 3779, 3782.5, 3786, 3789.5, 
    3793, 3796.5, 3800, 3803.5, 3807, 3810.5, 3814, 3817.4, 3820.9, 3824.4, 
    3827.9, 3831.3, 3834.8, 3838.3, 3841.8, 3845.2, 3848.7, 3852.2, 3855.7, 
    3859.1, 3862.6, 3866.1, 3869.5, 3873, 3876.5, 3879.9, 3883.4, 3886.8, 
    3890.3, 3893.7, 3897.2, 3900.6, 3904, 3907.4, 3910.8, 3914.2, 3917.7, 
    3921.1, 3924.5, 3927.9, 3931.3, 3934.7, 3938.2, 3941.6, 3945, 3948.4, 
    3951.9, 3955.3, 3958.7, 3962.1, 3965.6, 3969, 3972.4, 3975.8, 3979.3, 
    3982.7, 3986.1, 3989.5, 3992.9, 3996.3, 3999.7, 4003.1, 4006.6, 4010, 
    4013.4, 4016.8, 4020.2, 4023.7, 4027.1, 4030.5, 4033.9, 4037.4, 4040.8, 
    4044.3, 4047.7, 4051.1, 4054.6, 4058, 4061.5, 4064.9, 4068.4, 4071.8, 
    4075.3, 4078.8, 4082.2, 4085.7, 4089.2, 4092.7, 4096.1, 4099.6, 4103.1, 
    4106.6, 4110, 4113.5, 4117, 4120.5, 4123.9, 4127.4, 4130.9, 4134.4, 
    4137.9, 4141.3, 4144.8, 4148.3, 4151.7, 4155.2, 4158.7, 4162.2, 4165.6, 
    4169.1, 4172.5, 4176, 4179.5, 4182.9, 4186.4, 4189.8, 4193.3, 4196.7, 
    4200.1, 4203.6, 4207, 4210.4, 4213.8, 4217.2, 4220.6, 4224, 4227.4, 
    4230.8, 4234.2, 4237.6, 4241, 4244.4, 4247.8, 4251.2, 4254.6, 4258, 
    4261.4, 4264.8, 4268.2, 4271.6, 4275, 4278.3, 4281.7, 4285.1, 4288.5, 
    4291.9, 4295.2, 4298.6, 4302, 4305.4, 4308.8, 4312.1, 4315.5, 4318.9, 
    4322.3, 4325.7, 4329.1, 4332.5, 4335.8, 4339.2, 4342.6, 4346, 4349.4, 
    4352.9, 4356.3, 4359.7, 4363.1, 4366.5, 4370, 4373.4, 4376.8, 4380.2, 
    4383.6, 4387.1, 4390.5, 4393.9, 4397.3, 4400.8, 4404.2, 4407.6, 4411, 
    4414.4, 4417.9, 4421.3, 4424.7, 4428.1, 4431.6, 4435, 4438.4, 4441.8, 
    4445.3, 4448.7, 4452.1, 4455.6, 4459, 4462.4, 4465.9, 4469.3, 4472.8, 
    4476.2, 4479.6, 4483.1, 4486.5, 4490, 4493.4, 4496.8, 4500.2, 4503.7, 
    4507.1, 4510.5, 4513.9, 4517.3, 4520.7, 4524.1, 4527.6, 4531, 4534.4, 
    4537.8, 4541.2, 4544.6, 4548, 4551.4, 4554.8, 4558.2, 4561.6, 4565.1, 
    4568.5, 4571.9, 4575.3, 4578.7, 4582.1, 4585.4, 4588.8, 4592.2, 4595.6, 
    4599, 4602.3, 4605.7, 4609.1, 4612.4, 4615.8, 4619.1, 4622.5, 4625.9, 
    4629.2, 4632.6, 4636, 4639.4, 4642.7, 4646.1, 4649.5, 4652.9, 4656.3, 
    4659.7, 4663.1, 4666.5, 4669.8, 4673.2, 4676.6, 4680, 4683.5, 4686.9, 
    4690.3, 4693.7, 4697.1, 4700.6, 4704, 4707.4, 4710.8, 4714.3, 4717.7, 
    4721.1, 4724.6, 4728, 4731.4, 4734.9, 4738.3, 4741.7, 4745.2, 4748.6, 
    4752, 4755.5, 4758.9, 4762.3, 4765.8, 4769.2, 4772.7, 4776.1, 4779.5, 
    4783, 4786.4, 4789.9, 4793.3, 4796.7, 4800.2, 4803.6, 4807, 4810.5, 
    4813.9, 4817.3, 4820.8, 4824.2, 4827.6, 4831, 4834.4, 4837.8, 4841.3, 
    4844.7, 4848.1, 4851.5, 4855, 4858.4, 4861.8, 4865.3, 4868.7, 4872.1, 
    4875.6, 4879, 4882.4, 4885.8, 4889.2, 4892.7, 4896.1, 4899.5, 4902.9, 
    4906.3, 4909.7, 4913.1, 4916.5, 4920, 4923.4, 4926.8, 4930.2, 4933.6, 
    4937, 4940.4, 4943.8, 4947.3, 4950.7, 4954.1, 4957.5, 4960.9, 4964.4, 
    4967.8, 4971.2, 4974.6, 4978, 4981.5, 4984.9, 4988.3, 4991.7, 4995.1, 
    4998.5, 5001.9, 5005.4, 5008.8, 5012.2, 5015.6, 5019.1, 5022.5, 5025.9, 
    5029.4, 5032.8, 5036.2, 5039.7, 5043.1, 5046.5, 5049.9, 5053.4, 5056.8, 
    5060.2, 5063.7, 5067.1, 5070.5, 5074, 5077.4, 5080.9, 5084.3, 5087.8, 
    5091.2, 5094.6, 5098, 5101.5, 5104.9, 5108.3, 5111.7, 5115.1, 5118.6, 
    5122, 5125.4, 5128.8, 5132.2, 5135.6, 5139, 5142.4, 5145.8, 5149.2, 
    5152.6, 5156, 5159.4, 5162.8, 5166.2, 5169.6, 5172.9, 5176.3, 5179.7, 
    5183.1, 5186.4, 5189.8, 5193.2, 5196.5, 5199.9, 5203.2, 5206.6, 5209.9, 
    5213.3, 5216.6, 5220, 5223.4, 5226.7, 5230.1, 5233.4, 5236.8, 5240.1, 
    5243.5, 5246.8, 5250.2, 5253.6, 5256.9, 5260.3, 5263.6, 5267, 5270.3, 
    5273.7, 5277.1, 5280.4, 5283.8, 5287.2, 5290.5, 5293.9, 5297.3, 5300.6, 
    5304, 5307.4, 5310.7, 5314.1, 5317.5, 5320.9, 5324.3, 5327.6, 5331, 
    5334.4, 5337.8, 5341.1, 5344.5, 5347.9, 5351.3, 5354.6, 5358, 5361.4, 
    5364.8, 5368.1, 5371.5, 5374.9, 5378.2, 5381.6, 5385, 5388.3, 5391.7, 
    5395.1, 5398.5, 5401.8, 5405.2, 5408.5, 5411.9, 5415.3, 5418.6, 5422, 
    5425.4, 5428.7, 5432.1, 5435.4, 5438.8, 5442.2, 5445.5, 5448.9, 5452.3, 
    5455.6, 5459, 5462.4, 5465.7, 5469.1, 5472.5, 5475.8, 5479.2, 5482.6, 
    5486, 5489.3, 5492.7, 5496.1, 5499.5, 5502.9, 5506.2, 5509.6, 5513, 
    5516.4, 5519.8, 5523.2, 5526.5, 5529.9, 5533.3, 5536.7, 5540.1, 5543.5, 
    5546.8, 5550.2, 5553.6, 5557, 5560.4, 5563.7, 5567.1, 5570.5, 5573.9, 
    5577.2, 5580.6, 5584, 5587.3, 5590.7, 5594, 5597.4, 5600.8, 5604.1, 
    5607.5, 5610.8, 5614.2, 5617.5, 5620.9, 5624.3, 5627.6, 5631, 5634.3, 
    5637.7, 5641.1, 5644.4, 5647.8, 5651.1, 5654.5, 5657.8, 5661.2, 5664.5, 
    5667.9, 5671.2, 5674.5, 5677.9, 5681.2, 5684.6, 5687.9, 5691.3, 5694.6, 
    5698, 5701.3, 5704.7, 5708, 5711.4, 5714.7, 5718.1, 5721.4, 5724.8, 
    5728.1, 5731.5, 5734.9, 5738.2, 5741.6, 5744.9, 5748.2, 5751.6, 5754.9, 
    5758.3, 5761.6, 5765, 5768.3, 5771.6, 5775, 5778.3, 5781.7, 5785, 5788.4, 
    5791.7, 5795.1, 5798.4, 5801.8, 5805.1, 5808.5, 5811.8, 5815.2, 5818.5, 
    5821.9, 5825.2, 5828.6, 5831.9, 5835.3, 5838.6, 5842, 5845.4, 5848.7, 
    5852.1, 5855.4, 5858.7, 5862.1, 5865.4, 5868.8, 5872.1, 5875.5, 5878.8, 
    5882.2, 5885.5, 5888.9, 5892.2, 5895.6, 5898.9, 5902.2, 5905.6, 5908.9, 
    5912.3, 5915.7, 5919, 5922.4, 5925.7, 5929.1, 5932.4, 5935.8, 5939.2, 
    5942.5, 5945.9, 5949.3, 5952.7, 5956, 5959.4, 5962.8, 5966.1, 5969.5, 
    5972.9, 5976.3, 5979.7, 5983, 5986.4, 5989.8, 5993.2, 5996.6, 5999.9, 
    6003.3, 6006.7, 6010.1, 6013.5, 6016.8, 6020.2, 6023.6, 6027, 6030.4, 
    6033.7, 6037.1, 6040.5, 6043.9, 6047.3, 6050.7, 6054.1, 6057.4, 6060.8, 
    6064.2, 6067.6, 6071, 6074.3, 6077.7, 6081.1, 6084.5, 6087.8, 6091.2, 
    6094.6, 6097.9, 6101.3, 6104.6, 6108, 6111.3, 6114.7, 6118, 6121.4, 
    6124.8, 6128.1, 6131.5, 6134.9, 6138.2, 6141.6, 6144.9, 6148.3, 6151.6, 
    6155, 6158.3, 6161.7, 6165, 6168.4, 6171.7, 6175, 6178.4, 6181.7, 6185, 
    6188.4, 6191.7, 6195, 6198.3, 6201.7, 6205, 6208.3, 6211.7, 6215, 6218.3, 
    6221.7, 6225, 6228.4, 6231.7, 6235.1, 6238.4, 6241.7, 6245.1, 6248.4, 
    6251.8, 6255.1, 6258.4, 6261.8, 6265.1, 6268.4, 6271.8, 6275.1, 6278.4, 
    6281.8, 6285.1, 6288.5, 6291.8, 6295.1, 6298.5, 6301.8, 6305.2, 6308.5, 
    6311.9, 6315.2, 6318.6, 6321.9, 6325.3, 6328.6, 6332, 6335.4, 6338.7, 
    6342.1, 6345.4, 6348.8, 6352.1, 6355.4, 6358.8, 6362.1, 6365.5, 6368.8, 
    6372.2, 6375.5, 6378.9, 6382.2, 6385.6, 6389, 6392.4, 6395.7, 6399.1, 
    6402.5, 6405.8, 6409.2, 6412.5, 6415.9, 6419.3, 6422.7, 6426, 6429.4, 
    6432.8, 6436.1, 6439.5, 6442.9, 6446.3, 6449.6, 6453, 6456.4, 6459.8, 
    6463.1, 6466.5, 6469.9, 6473.3, 6476.6, 6480, 6483.4, 6486.8, 6490.1, 
    6493.5, 6496.9, 6500.3, 6503.6, 6507, 6510.4, 6513.8, 6517.1, 6520.5, 
    6523.9, 6527.2, 6530.6, 6534, 6537.4, 6540.7, 6544.1, 6547.5, 6550.8, 
    6554.2, 6557.5, 6560.8, 6564.2, 6567.5, 6570.9, 6574.2, 6577.5, 6580.9, 
    6584.2, 6587.5, 6590.8, 6594.2, 6597.5, 6600.8, 6604.1, 6607.4, 6610.8, 
    6614.1, 6617.4, 6620.7, 6624, 6627.3, 6630.6, 6633.9, 6637.2, 6640.5, 
    6643.8, 6647.1, 6650.4, 6653.7, 6656.9, 6660.2, 6663.5, 6666.8, 6670, 
    6673.3, 6676.6, 6679.9, 6683.1, 6686.4, 6689.7, 6693, 6696.3, 6699.5, 
    6702.8, 6706.1, 6709.4, 6712.7, 6716, 6719.2, 6722.5, 6725.8, 6729.1, 
    6732.4, 6735.7, 6738.9, 6742.2, 6745.5, 6748.8, 6752.1, 6755.4, 6758.7, 
    6762, 6765.3, 6768.6, 6771.9, 6775.2, 6778.5, 6781.8, 6785.1, 6788.4, 
    6791.7, 6795.1, 6798.4, 6801.7, 6805, 6808.3, 6811.6, 6814.9, 6818.2, 
    6821.6, 6824.9, 6828.2, 6831.5, 6834.8, 6838.1, 6841.5, 6844.8, 6848.1, 
    6851.4, 6854.7, 6858.1, 6861.4, 6864.7, 6868, 6871.4, 6874.7, 6878, 
    6881.4, 6884.7, 6888, 6891.4, 6894.7, 6898, 6901.4, 6904.7, 6908, 6911.4, 
    6914.7, 6918, 6921.4, 6924.7, 6928, 6931.4, 6934.7, 6938.1, 6941.4, 
    6944.7, 6948.1, 6951.4, 6954.8, 6958.1, 6961.5, 6964.8, 6968.2, 6971.5, 
    6974.9, 6978.2, 6981.6, 6984.9, 6988.2, 6991.6, 6994.9, 6998.3, 7001.6, 
    7005, 7008.3, 7011.6, 7015, 7018.3, 7021.7, 7025, 7028.4, 7031.7, 7035, 
    7038.4, 7041.7, 7045.1, 7048.4, 7051.8, 7055.1, 7058.5, 7061.8, 7065.2, 
    7068.5, 7071.9, 7075.2, 7078.5, 7081.9, 7085.2, 7088.5, 7091.9, 7095.2, 
    7098.5, 7101.8, 7105.2, 7108.5, 7111.8, 7115.2, 7118.5, 7121.8, 7125.2, 
    7128.5, 7131.8, 7135.2, 7138.5, 7141.8, 7145.2, 7148.5, 7151.8, 7155.2, 
    7158.5, 7161.8, 7165.2, 7168.5, 7171.8, 7175.1, 7178.4, 7181.8, 7185.1, 
    7188.4, 7191.7, 7195, 7198.4, 7201.7, 7205, 7208.3, 7211.7, 7215, 7218.3, 
    7221.6, 7225, 7228.3, 7231.7, 7235, 7238.3, 7241.7, 7245, 7248.3, 7251.7, 
    7255, 7258.4, 7261.7, 7265, 7268.4, 7271.7, 7275, 7278.3, 7281.7, 7285, 
    7288.3, 7291.6, 7295, 7298.3, 7301.6, 7304.9, 7308.3, 7311.6, 7314.9, 
    7318.3, 7321.6, 7324.9, 7328.3, 7331.6, 7334.9, 7338.3, 7341.6, 7344.9, 
    7348.2, 7351.5, 7354.9, 7358.2, 7361.5, 7364.8, 7368.1, 7371.4, 7374.8, 
    7378.1, 7381.4, 7384.7, 7388, 7391.3, 7394.6, 7397.9, 7401.2, 7404.5, 
    7407.9, 7411.2, 7414.5, 7417.8, 7421.1, 7424.4, 7427.7, 7431.1, 7434.4, 
    7437.7, 7441, 7444.3, 7447.6, 7450.9, 7454.2, 7457.5, 7460.8, 7464.1, 
    7467.4, 7470.7, 7474, 7477.3, 7480.6, 7483.9, 7487.3, 7490.6, 7493.9, 
    7497.2, 7500.5, 7503.8, 7507.1, 7510.4, 7513.7, 7517, 7520.3, 7523.6, 
    7526.9, 7530.2, 7533.5, 7536.8, 7540.1, 7543.4, 7546.7, 7550, 7553.3, 
    7556.6, 7559.9, 7563.2, 7566.5, 7569.8, 7573.1, 7576.5, 7579.8, 7583.1, 
    7586.4, 7589.7, 7593, 7596.4, 7599.7, 7603, 7606.3, 7609.6, 7612.9, 
    7616.2, 7619.6, 7622.9, 7626.2, 7629.5, 7632.8, 7636.1, 7639.4, 7642.7, 
    7646, 7649.4, 7652.7, 7656, 7659.3, 7662.6, 7665.9, 7669.2, 7672.6, 
    7675.9, 7679.2, 7682.5, 7685.8, 7689.1, 7692.5, 7695.8, 7699.1, 7702.4, 
    7705.7, 7709, 7712.3, 7715.6, 7718.9, 7722.2, 7725.5, 7728.8, 7732.1, 
    7735.4, 7738.7, 7742, 7745.3, 7748.6, 7751.9, 7755.2, 7758.5, 7761.8, 
    7765.1, 7768.4, 7771.7, 7775, 7778.3, 7781.6, 7784.9, 7788.2, 7791.5, 
    7794.8, 7798.1, 7801.4, 7804.7, 7808, 7811.3, 7814.6, 7817.9, 7821.2, 
    7824.4, 7827.7, 7831, 7834.3, 7837.5, 7840.8, 7844.1, 7847.4, 7850.7, 
    7854, 7857.3, 7860.6, 7863.8, 7867.1, 7870.4, 7873.7, 7877, 7880.3, 
    7883.6, 7886.9, 7890.2, 7893.4, 7896.7, 7900, 7903.3, 7906.5, 7909.8, 
    7913.1, 7916.4, 7919.6, 7922.9, 7926.2, 7929.4, 7932.7, 7936, 7939.2, 
    7942.5, 7945.8, 7949.1, 7952.3, 7955.6, 7958.9, 7962.2, 7965.4, 7968.7, 
    7972, 7975.3, 7978.5, 7981.8, 7985.1, 7988.4, 7991.6, 7994.9, 7998.2, 
    8001.5, 8004.7, 8008, 8011.3, 8014.6, 8017.9, 8021.2, 8024.5, 8027.7, 
    8031, 8034.3, 8037.6, 8040.9, 8044.2, 8047.5, 8050.9, 8054.2, 8057.4, 
    8060.7, 8064, 8067.3, 8070.6, 8073.9, 8077.2, 8080.5, 8083.7, 8087, 
    8090.3, 8093.6, 8096.9, 8100.2, 8103.4, 8106.7, 8110, 8113.3, 8116.6, 
    8119.8, 8123.1, 8126.4, 8129.7, 8132.9, 8136.2, 8139.5, 8142.8, 8146, 
    8149.3, 8152.6, 8155.8, 8159.1, 8162.4, 8165.6, 8168.9, 8172.1, 8175.4, 
    8178.6, 8181.9, 8185.2, 8188.4, 8191.7, 8194.9, 8198.2, 8201.4, 8204.7, 
    8207.9, 8211.2, 8214.5, 8217.8, 8221, 8224.3, 8227.6, 8230.8, 8234.1, 
    8237.4, 8240.7, 8243.9, 8247.2, 8250.5, 8253.8, 8257.1, 8260.3, 8263.6, 
    8266.9, 8270.2, 8273.4, 8276.7, 8280, 8283.3, 8286.6, 8289.9, 8293.1, 
    8296.4, 8299.7, 8303, 8306.3, 8309.6, 8312.9, 8316.2, 8319.5, 8322.8, 
    8326.1, 8329.4, 8332.6, 8335.9, 8339.2, 8342.5, 8345.8, 8349.1, 8352.4, 
    8355.7, 8359, 8362.3, 8365.6, 8368.9, 8372.2, 8375.5, 8378.8, 8382.1, 
    8385.3, 8388.6, 8391.9, 8395.2, 8398.5, 8401.8, 8405, 8408.3, 8411.6, 
    8414.9, 8418.1, 8421.4, 8424.7, 8428, 8431.3, 8434.5, 8437.8, 8441.1, 
    8444.4, 8447.6, 8450.9, 8454.2, 8457.5, 8460.7, 8464, 8467.3, 8470.6, 
    8473.9, 8477.1, 8480.4, 8483.7, 8486.9, 8490.2, 8493.5, 8496.7, 8500, 
    8503.3, 8506.5, 8509.8, 8513.1, 8516.3, 8519.6, 8522.9, 8526.2, 8529.4, 
    8532.7, 8536, 8539.2, 8542.5, 8545.8, 8549, 8552.3, 8555.5, 8558.8, 
    8562.1, 8565.3, 8568.6, 8571.9, 8575.1, 8578.4, 8581.7, 8584.9, 8588.2, 
    8591.4, 8594.7, 8598, 8601.2, 8604.5, 8607.7, 8611, 8614.3, 8617.5, 
    8620.8, 8624.1, 8627.4, 8630.7, 8633.9, 8637.2, 8640.5, 8643.8, 8647.1, 
    8650.4, 8653.6, 8656.9, 8660.2, 8663.5, 8666.8, 8670.1, 8673.3, 8676.6, 
    8679.9, 8683.2, 8686.5, 8689.8, 8693.1, 8696.4, 8699.7, 8702.9, 8706.2, 
    8709.5, 8712.8, 8716.1, 8719.4, 8722.7, 8726, 8729.3, 8732.6, 8735.9, 
    8739.2, 8742.5, 8745.8, 8749.1, 8752.4, 8755.7, 8758.9, 8762.2, 8765.5, 
    8768.8, 8772.1, 8775.3, 8778.6, 8781.9, 8785.2, 8788.5, 8791.8, 8795, 
    8798.3, 8801.6, 8804.9, 8808.2, 8811.5, 8814.8, 8818.1, 8821.4, 8824.6, 
    8827.9, 8831.2, 8834.5, 8837.7, 8841, 8844.3, 8847.5, 8850.8, 8854, 
    8857.3, 8860.5, 8863.8, 8867, 8870.3, 8873.5, 8876.8, 8880, 8883.3, 
    8886.6, 8889.8, 8893.1, 8896.3, 8899.6, 8902.8, 8906.1, 8909.3, 8912.6, 
    8915.8, 8919.1, 8922.3, 8925.5, 8928.8, 8932, 8935.3, 8938.5, 8941.7, 
    8945, 8948.2, 8951.5, 8954.7, 8958, 8961.2, 8964.5, 8967.7, 8971, 8974.2, 
    8977.5, 8980.7, 8984, 8987.2, 8990.4, 8993.7, 8996.9, 9000.2, 9003.4, 
    9006.6, 9009.9, 9013.1, 9016.3, 9019.6, 9022.8, 9026, 9029.3, 9032.5, 
    9035.8, 9039, 9042.2, 9045.5, 9048.7, 9052, 9055.2, 9058.4, 9061.7, 
    9064.9, 9068.2, 9071.4, 9074.6, 9077.9, 9081.1, 9084.3, 9087.6, 9090.8, 
    9094.1, 9097.3, 9100.6, 9103.8, 9107, 9110.3, 9113.5, 9116.8, 9120, 
    9123.3, 9126.5, 9129.8, 9133, 9136.3, 9139.5, 9142.8, 9146, 9149.3, 
    9152.5, 9155.8, 9159, 9162.3, 9165.5, 9168.8, 9172, 9175.3, 9178.5, 
    9181.8, 9185.1, 9188.3, 9191.6, 9194.8, 9198.1, 9201.3, 9204.6, 9207.8, 
    9211.1, 9214.3, 9217.6, 9220.8, 9224.1, 9227.3, 9230.6, 9233.9, 9237.1, 
    9240.4, 9243.7, 9246.9, 9250.2, 9253.5, 9256.7, 9260, 9263.2, 9266.5, 
    9269.8, 9273, 9276.3, 9279.6, 9282.9, 9286.1, 9289.4, 9292.7, 9295.9, 
    9299.2, 9302.5, 9305.8, 9309, 9312.3, 9315.5, 9318.8, 9322.1, 9325.3, 
    9328.6, 9331.9, 9335.1, 9338.4, 9341.6, 9344.9, 9348.1, 9351.4, 9354.7, 
    9357.9, 9361.2, 9364.4, 9367.7, 9370.9, 9374.2, 9377.5, 9380.7, 9384, 
    9387.2, 9390.5, 9393.7, 9397, 9400.2, 9403.5, 9406.7, 9410, 9413.2, 
    9416.5, 9419.7, 9423, 9426.3, 9429.5, 9432.8, 9436, 9439.3, 9442.5, 
    9445.8, 9449.1, 9452.3, 9455.6, 9458.9, 9462.1, 9465.4, 9468.6, 9471.9, 
    9475.2, 9478.4, 9481.7, 9485, 9488.2, 9491.5, 9494.7, 9498, 9501.3, 
    9504.5, 9507.8, 9511, 9514.3, 9517.6, 9520.8, 9524.1, 9527.3, 9530.6, 
    9533.9, 9537.1, 9540.4, 9543.7, 9546.9, 9550.2, 9553.4, 9556.7, 9560, 
    9563.2, 9566.5, 9569.8, 9573, 9576.3, 9579.5, 9582.8, 9586.1, 9589.3, 
    9592.6, 9595.9, 9599.1, 9602.4, 9605.7, 9608.9, 9612.2, 9615.5, 9618.8, 
    9622, 9625.3, 9628.6, 9631.8, 9635.1, 9638.3, 9641.6, 9644.9, 9648.1, 
    9651.4, 9654.6, 9657.9, 9661.1, 9664.3, 9667.6, 9670.8, 9674.1, 9677.3, 
    9680.6, 9683.8, 9687.1, 9690.3, 9693.6, 9696.8, 9700.1, 9703.3, 9706.6, 
    9709.8, 9713.1, 9716.3, 9719.6, 9722.8, 9726.1, 9729.3, 9732.6, 9735.8, 
    9739, 9742.3, 9745.5, 9748.8, 9752, 9755.2, 9758.5, 9761.7, 9764.9, 
    9768.2, 9771.4, 9774.7, 9777.9, 9781.1, 9784.4, 9787.6, 9790.9, 9794.1, 
    9797.4, 9800.6, 9803.8, 9807.1, 9810.3, 9813.5, 9816.8, 9820, 9823.2, 
    9826.5, 9829.7, 9832.9, 9836.2, 9839.4, 9842.6, 9845.9, 9849.1, 9852.4, 
    9855.6, 9858.8, 9862.1, 9865.3, 9868.5, 9871.7, 9875, 9878.2, 9881.4, 
    9884.7, 9887.9, 9891.2, 9894.4, 9897.6, 9900.9, 9904.1, 9907.4, 9910.6, 
    9913.8, 9917.1, 9920.3, 9923.6, 9926.8, 9930.1, 9933.3, 9936.5, 9939.8, 
    9943, 9946.2, 9949.5, 9952.7, 9955.9, 9959.2, 9962.4, 9965.6, 9968.9, 
    9972.1, 9975.4, 9978.6, 9981.8, 9985.1, 9988.3, 9991.6, 9994.8, 9998.1, 
    10001, 10005, 10008, 10011, 10014, 10018, 10021, 10024, 10027, 10031, 
    10034, 10037, 10040, 10043, 10047, 10050, 10053, 10056, 10060, 10063, 
    10066, 10069, 10073, 10076, 10079, 10082, 10086, 10089, 10092, 10095, 
    10098, 10102, 10105, 10108, 10111, 10115, 10118, 10121, 10124, 10128, 
    10131, 10134, 10137, 10140, 10144, 10147, 10150, 10153, 10157, 10160, 
    10163, 10166, 10170, 10173, 10176, 10179, 10183, 10186, 10189, 10192, 
    10195, 10199, 10202, 10205, 10208, 10212, 10215, 10218, 10221, 10225, 
    10228, 10231, 10234, 10238, 10241, 10244, 10247, 10250, 10254, 10257, 
    10260, 10263, 10267, 10270, 10273, 10276, 10279, 10283, 10286, 10289, 
    10292, 10296, 10299, 10302, 10305, 10308, 10312, 10315, 10318, 10321, 
    10324, 10328, 10331, 10334, 10337, 10340, 10344, 10347, 10350, 10353, 
    10357, 10360, 10363, 10366, 10369, 10373, 10376, 10379, 10382, 10386, 
    10389, 10392, 10395, 10399, 10402, 10405, 10408, 10411, 10415, 10418, 
    10421, 10424, 10428, 10431, 10434, 10437, 10441, 10444, 10447, 10450, 
    10454, 10457, 10460, 10463, 10467, 10470, 10473, 10476, 10480, 10483, 
    10486, 10489, 10493, 10496, 10499, 10503, 10506, 10509, 10512, 10516, 
    10519, 10522, 10525, 10529, 10532, 10535, 10538, 10542, 10545, 10548, 
    10552, 10555, 10558, 10561, 10565, 10568, 10571, 10575, 10578, 10581, 
    10584, 10588, 10591, 10594, 10597, 10601, 10604, 10607, 10611, 10614, 
    10617, 10620, 10624, 10627, 10630, 10634, 10637, 10640, 10643, 10647, 
    10650, 10653, 10657, 10660, 10663, 10666, 10670, 10673, 10676, 10680, 
    10683, 10686, 10689, 10693, 10696, 10699, 10703, 10706, 10709, 10712, 
    10716, 10719, 10722, 10726, 10729, 10732, 10736, 10739, 10742, 10745, 
    10749, 10752, 10755, 10759, 10762, 10765, 10769, 10772, 10775, 10778, 
    10782, 10785, 10788, 10792, 10795, 10798, 10802, 10805, 10808, 10812, 
    10815, 10818, 10822, 10825, 10828, 10831, 10835, 10838, 10841, 10845, 
    10848, 10851, 10855, 10858, 10861, 10865, 10868, 10871, 10875, 10878, 
    10881, 10885, 10888, 10891, 10894, 10898, 10901, 10904, 10908, 10911, 
    10914, 10918, 10921, 10924, 10928, 10931, 10934, 10938, 10941, 10944, 
    10948, 10951, 10954, 10958, 10961, 10964, 10968, 10971, 10974, 10978, 
    10981, 10984, 10988, 10991, 10994, 10997, 11001, 11004, 11007, 11011, 
    11014, 11017, 11020, 11024, 11027, 11030, 11033, 11037, 11040, 11043, 
    11046, 11050, 11053, 11056, 11059, 11063, 11066, 11069, 11072, 11075, 
    11079, 11082, 11085, 11088, 11091, 11095, 11098, 11101, 11104, 11107, 
    11111, 11114, 11117, 11120, 11124, 11127, 11130, 11133, 11136, 11140, 
    11143, 11146, 11149, 11153, 11156, 11159, 11162, 11165, 11169, 11172, 
    11175, 11178, 11182, 11185, 11188, 11191, 11194, 11198, 11201, 11204, 
    11207, 11210, 11214, 11217, 11220, 11223, 11227, 11230, 11233, 11236, 
    11239, 11243, 11246, 11249, 11252, 11255, 11259, 11262, 11265, 11268, 
    11271, 11275, 11278, 11281, 11284, 11287, 11291, 11294, 11297, 11300, 
    11304, 11307, 11310, 11313, 11316, 11320, 11323, 11326, 11329, 11333, 
    11336, 11339, 11342, 11346, 11349, 11352, 11355, 11359, 11362, 11365, 
    11368, 11372, 11375, 11378, 11382, 11385, 11388, 11391, 11395, 11398, 
    11401, 11405, 11408, 11411, 11414, 11418, 11421, 11424, 11427, 11431, 
    11434, 11437, 11441, 11444, 11447, 11450, 11454, 11457, 11460, 11463, 
    11467, 11470, 11473, 11477, 11480, 11483, 11486, 11490, 11493, 11496, 
    11499, 11503, 11506, 11509, 11512, 11516, 11519, 11522, 11525, 11529, 
    11532, 11535, 11539, 11542, 11545, 11548, 11552, 11555, 11558, 11562, 
    11565, 11568, 11571, 11575, 11578, 11581, 11585, 11588, 11591, 11594, 
    11598, 11601, 11604, 11607, 11611, 11614, 11617, 11621, 11624, 11627, 
    11630, 11634, 11637, 11640, 11643, 11647, 11650, 11653, 11656, 11660, 
    11663, 11666, 11669, 11672, 11676, 11679, 11682, 11685, 11689, 11692, 
    11695, 11698, 11702, 11705, 11708, 11711, 11715, 11718, 11721, 11725, 
    11728, 11731, 11734, 11738, 11741, 11744, 11748, 11751, 11754, 11757, 
    11761, 11764, 11767, 11770, 11774, 11777, 11780, 11784, 11787, 11790, 
    11793, 11797, 11800, 11803, 11807, 11810, 11813, 11816, 11820, 11823, 
    11826, 11829, 11833, 11836, 11839, 11842, 11846, 11849, 11852, 11855, 
    11859, 11862, 11865, 11869, 11872, 11875, 11878, 11882, 11885, 11888, 
    11891, 11895, 11898, 11901, 11904, 11908, 11911, 11914, 11918, 11921, 
    11924, 11927, 11931, 11934, 11937, 11941, 11944, 11947, 11950, 11954, 
    11957, 11960, 11963, 11967, 11970, 11973, 11976, 11980, 11983, 11986, 
    11989, 11993, 11996, 11999, 12002, 12006, 12009, 12012, 12015, 12019, 
    12022, 12025, 12028, 12032, 12035, 12038, 12041, 12045, 12048, 12051, 
    12054, 12058, 12061, 12064, 12067, 12071, 12074, 12077, 12080, 12084, 
    12087, 12090, 12093, 12096, 12100, 12103, 12106, 12109, 12113, 12116, 
    12119, 12122, 12125, 12129, 12132, 12135, 12138, 12141, 12145, 12148, 
    12151, 12154, 12157, 12161, 12164, 12167, 12170, 12173, 12177, 12180, 
    12183, 12186, 12189, 12193, 12196, 12199, 12202, 12205, 12209, 12212, 
    12215, 12218, 12221, 12225, 12228, 12231, 12234, 12238, 12241, 12244, 
    12247, 12250, 12254, 12257, 12260, 12263, 12267, 12270, 12273, 12276, 
    12280, 12283, 12286, 12289, 12292, 12296, 12299, 12302, 12305, 12309, 
    12312, 12315, 12318, 12322, 12325, 12328, 12331, 12335, 12338, 12341, 
    12344, 12347, 12351, 12354, 12357, 12360, 12364, 12367, 12370, 12373, 
    12376, 12380, 12383, 12386, 12389, 12393, 12396, 12399, 12402, 12406, 
    12409, 12412, 12415, 12419, 12422, 12425, 12428, 12431, 12435, 12438, 
    12441, 12444, 12448, 12451, 12454, 12457, 12461, 12464, 12467, 12470, 
    12473, 12477, 12480, 12483, 12486, 12489, 12493, 12496, 12499, 12502, 
    12505, 12509, 12512, 12515, 12518, 12521, 12525, 12528, 12531, 12534, 
    12537, 12541, 12544, 12547, 12550, 12553, 12557, 12560, 12563, 12566, 
    12569, 12573, 12576, 12579, 12582, 12585, 12589, 12592, 12595, 12598, 
    12601, 12605, 12608, 12611, 12614, 12617, 12621, 12624, 12627, 12630, 
    12633, 12637, 12640, 12643, 12646, 12650, 12653, 12656, 12659, 12662, 
    12666, 12669, 12672, 12675, 12678, 12682, 12685, 12688, 12691, 12694, 
    12698, 12701, 12704, 12707, 12711, 12714, 12717, 12720, 12723, 12727, 
    12730, 12733, 12736, 12739, 12743, 12746, 12749, 12752, 12755, 12759, 
    12762, 12765, 12768, 12771, 12775, 12778, 12781, 12784, 12787, 12791, 
    12794, 12797, 12800, 12803, 12806, 12810, 12813, 12816, 12819, 12822, 
    12825, 12829, 12832, 12835, 12838, 12841, 12845, 12848, 12851, 12854, 
    12857, 12860, 12864, 12867, 12870, 12873, 12876, 12879, 12883, 12886, 
    12896, 12907, 12917, 12927, 12937, 12947, 12957, 12966, 12976, 12985, 
    12995, 13004, 13014, 13024, 13034, 13044, 13055, 13066, 13077, 13088, 
    13100, 13112, 13124, 13136, 13149, 13162, 13175, 13188, 13201, 13214, 
    13228, 13241, 13254, 13267, 13280, 13292, 13305, 13317, 13329, 13341, 
    13353, 13365, 13377, 13388, 13400, 13411, 13423, 13434, 13446, 13457, 
    13469, 13480, 13492, 13504, 13516, 13528, 13540, 13552, 13565, 13577, 
    13590, 13602, 13615, 13628, 13640, 13653, 13666, 13679, 13691, 13704, 
    13717, 13729, 13742, 13754, 13767, 13779, 13791, 13803, 13816, 13828, 
    13840, 13852, 13864, 13877, 13889, 13901, 13914, 13926, 13939, 13951, 
    13964, 13977, 13990, 14003, 14016, 14029, 14043, 14056, 14069, 14083, 
    14096, 14110, 14123, 14137, 14150, 14164, 14178, 14191, 14205, 14218, 
    14232, 14246, 14259, 14273, 14286, 14300, 14313, 14327, 14340, 14354, 
    14367, 14380, 14394, 14407, 14420, 14433, 14446, 14460, 14473, 14486, 
    14499, 14512, 14525, 14538, 14551, 14564, 14577, 14590, 14603, 14616, 
    14629, 14642, 14656, 14669, 14683, 14696, 14710, 14724, 14738, 14752, 
    14766, 14780, 14795, 14810, 14824, 14839, 14854, 14870, 14885, 14900, 
    14916, 14931, 14947, 14962, 14978, 14994, 15010, 15025, 15041, 15057, 
    15073, 15089, 15104, 15120, 15136, 15152, 15167, 15183, 15199, 15214, 
    15230, 15246, 15261, 15277, 15293, 15308, 15324, 15339, 15355, 15371, 
    15386, 15402, 15418, 15433, 15449, 15464, 15480, 15496, 15512, 15527, 
    15543, 15559, 15575, 15591, 15607, 15624, 15640, 15657, 15674, 15691, 
    15709, 15727, 15745, 15763, 15781, 15800, 15819, 15838, 15858, 15878, 
    15898, 15918, 15938, 15958, 15979, 16000, 16020, 16041, 16062, 16082, 
    16103, 16124, 16145, 16165, 16186, 16207, 16227, 16248, 16268, 16289, 
    16309, 16329, 16350, 16370, 16390, 16410, 16431, 16451, 16471, 16490, 
    16510, 16530, 16549, 16568, 16588, 16607, 16625, 16644, 16662, 16680, 
    16698, 16715, 16732, 16749, 16766, 16783, 16799, 16815, 16831, 16847, 
    16862, 16877, 16893, 16908, 16923, 16938, 16953, 16968, 16983, 16998, 
    17013, 17028, 17043, 17059, 17074, 17089, 17105, 17120, 17136, 17151, 
    17167, 17183, 17198, 17214, 17229, 17245, 17261, 17277, 17292, 17308, 
    17324, 17341, 17357, 17373, 17390, 17407, 17424, 17441, 17459, 17476, 
    17494, 17512, 17531, 17550, 17569, 17588, 17607, 17627, 17647, 17667, 
    17687, 17707, 17728, 17749, 17770, 17791, 17813, 17835, 17856, 17878, 
    17900, 17922, 17945, 17967, 17990, 18012, 18035, 18057, 18080, 18103, 
    18126, 18148, 18171, 18194, 18216, 18239, 18261, 18284, 18306, 18328, 
    18351, 18373, 18395, 18416, 18438, 18460, 18481, 18503, 18524, 18545, 
    18566, 18587, 18608, 18629, 18650, 18670, 18690, 18711, 18731, 18751, 
    18771, 18791, 18811, 18831, 18850, 18870, 18890, 18909, 18929, 18948, 
    18968, 18987, 19007, 19026, 19045, 19065, 19084, 19103, 19123, 19142, 
    19161, 19180, 19200, 19219, 19238, 19257, 19277, 19296, 19315, 19335, 
    19354, 19374, 19394, 19413, 19433, 19454, 19474, 19494, 19515, 19536, 
    19557, 19578, 19600, 19621, 19643, 19665, 19687, 19709, 19731, 19753, 
    19775, 19797, 19820, 19842, 19864, 19886, 19908, 19930, 19952, 19974, 
    19995, 20017, 20039, 20060, 20082, 20103, 20125, 20146, 20168, 20190, 
    20211, 20233, 20255, 20276, 20298, 20320, 20342, 20364, 20386, 20409, 
    20431, 20453, 20475, 20498, 20520, 20543, 20565, 20588, 20610, 20633, 
    20656, 20679, 20702, 20726, 20749, 20773, 20797, 20821, 20846, 20870, 
    20895, 20920, 20945, 20970, 20996, 21022, 21047, 21073, 21099, 21125, 
    21152, 21178, 21204, 21230, 21256, 21282, 21308, 21334, 21360, 21385, 
    21411, 21436, 21461, 21486, 21511, 21535, 21560, 21584, 21607, 21631, 
    21654, 21678, 21701, 21723, 21746, 21769, 21791, 21813, 21836, 21858, 
    21880, 21902, 21925, 21947, 21970, 21992, 22015, 22038, 22062, 22085, 
    22109, 22133, 22158, 22182, 22207, 22233, 22259, 22284, 22311, 22337, 
    22364, 22391, 22418, 22445, 22473, 22500, 22528, 22556, 22584, 22611, 
    22639, 22667, 22695, 22723, 22751, 22778, 22806, 22834, 22861, 22889, 
    22916, 22944, 22971, 22999, 23026, 23053, 23081, 23108, 23136, 23163, 
    23190, 23217, 23245, 23272, 23299, 23326, 23353, 23379, 23406, 23432, 
    23459, 23485, 23511, 23536, 23562, 23587, 23613, 23638, 23663, 23688, 
    23713, 23738, 23763, 23787, 23812, 23837, 23862, 23887, 23912, 23938, 
    23963, 23989, 24015, 24041, 24067, 24093, 24120, 24147, 24174, 24201, 
    24228, 24256, 24284, 24312, 24341, 24369, 24398, 24427, 24456, 24486, 
    24515, 24545, 24575, 24605, 24635, 24666, 24696, 24726, 24757, 24787, 
    24818, 24848, 24879, 24909, 24940, 24970, 25000, 25031, 25061, 25091, 
    25121, 25151, 25182, 25212, 25242, 25271, 25301, 25331, 25361, 25391, 
    25420, 25450, 25480, 25509, 25539, 25568, 25597, 25627, 25656, 25685, 
    25715, 25744, 25773, 25802, 25832, 25861, 25890, 25919, 25949, 25978, 
    26007, 26036, 26065, 26094, 26123, 26152, 26181, 26209, 26238, 26266, 
    26294, 26323, 26351, 26379, 26407, 26435, 26463, 26491, 26519, 26547, 
    26576, 26605, 26633, 26662, 26691, 26721, 26750, 26780, 26810, 26840, 
    26871, 26902, 26933, 26964, 26995, 27027, 27059, 27091, 27124, 27156, 
    27189, 27222, 27255, 27288, 27322, 27355, 27389, 27423, 27456, 27490, 
    27523, 27557, 27590, 27624, 27657, 27691, 27724, 27757, 27790, 27823, 
    27855, 27888, 27921, 27953, 27985, 28018, 28050, 28082, 28114, 28146, 
    28178, 28210, 28242, 28274, 28306, 28337, 28369, 28401, 28433, 28465, 
    28496, 28528, 28560, 28592, 28624, 28655, 28687, 28719, 28751, 28783, 
    28815, 28846, 28878, 28910, 28942, 28974, 29006, 29037, 29069, 29101, 
    29133, 29165, 29196, 29228, 29260, 29291, 29323, 29354, 29386, 29417, 
    29448, 29480, 29511, 29542, 29574, 29605, 29636, 29667, 29698, 29729, 
    29760, 29792, 29823, 29854, 29886, 29918, 29949, 29981, 30013, 30046, 
    30078, 30111, 30143, 30176, 30209, 30243, 30276, 30310, 30343, 30377, 
    30411, 30445, 30479, 30514, 30548, 30582, 30617, 30651, 30685, 30720, 
    30754, 30788, 30822, 30857, 30891, 30925, 30959, 30993, 31027, 31061, 
    31095, 31129, 31163, 31197, 31231, 31265, 31298, 31332, 31366, 31400, 
    31434, 31468, 31502, 31536, 31570, 31604, 31638, 31672, 31706, 31741, 
    31775, 31810, 31844, 31879, 31914, 31948, 31983, 32018, 32053, 32088, 
    32123, 32158, 32193, 32228, 32262, 32297, 32332, 32367, 32402, 32437, 
    32471, 32506, 32541, 32576, 32611, 32645, 32680, 32715, 32750, 32785, 
    32820, 32855, 32890, 32925, 32960, 32996, 33031, 33066, 33101, 33137, 
    33172, 33207, 33243, 33278, 33313, 33349, 33384, 33419, 33455, 33490, 
    33525, 33560, 33595, 33630, 33665, 33700, 33735, 33770, 33805, 33840, 
    33874, 33909, 33944, 33978, 34013, 34048, 34082, 34117, 34151, 34186, 
    34221, 34255, 34290, 34324, 34359, 34394, 34428, 34463, 34498, 34532, 
    34567, 34602, 34637, 34671, 34706, 34741, 34776, 34811, 34846, 34882, 
    34917, 34952, 34988, 35023, 35059, 35094, 35130, 35166, 35201, 35237, 
    35273, 35309, 35344, 35380, 35416, 35451, 35487, 35522, 35557, 35593, 
    35628, 35663, 35698, 35734, 35769, 35804, 35839, 35874, 35910, 35945, 
    35980, 36016, 36051, 36087, 36123, 36158, 36194, 36230, 36266, 36302, 
    36338, 36374, 36411, 36447, 36483, 36519, 36555, 36592, 36628, 36664, 
    36700, 36736, 36772, 36808, 36844, 36880, 36916, 36951, 36987, 37022, 
    37058, 37093, 37129, 37164, 37199, 37234, 37269, 37304, 37339, 37374, 
    37409, 37444, 37479, 37513, 37548, 37583, 37618, 37653, 37688, 37723, 
    37758, 37794, 37829, 37864, 37900, 37935, 37971, 38007, 38043, 38079, 
    38115, 38151, 38187, 38224, 38260, 38297, 38334, 38370, 38407, 38444, 
    38481, 38518, 38555, 38592, 38629, 38666, 38703, 38740, 38776, 38813, 
    38850, 38887, 38924, 38960, 38997, 39034, 39070, 39107, 39143, 39180, 
    39216, 39252, 39288, 39325, 39361, 39397, 39433, 39469, 39506, 39542, 
    39578, 39614, 39650, 39686, 39722, 39757, 39793, 39829, 39865, 39901, 
    39937, 39973, 40008, 40044, 40080, 40116, 40152, 40188, 40224, 40260, 
    40296, 40331, 40367, 40403, 40439, 40475, 40511, 40548, 40584, 40620, 
    40656, 40692, 40728, 40764, 40800, 40836, 40872, 40909, 40945, 40981, 
    41017, 41053, 41090, 41126, 41162, 41199, 41235, 41271, 41308, 41344, 
    41381, 41417, 41454, 41490, 41527, 41563, 41599, 41636, 41672, 41709, 
    41745, 41782, 41818, 41855, 41891, 41928, 41964, 42000, 42037, 42073, 
    42110, 42146, 42182, 42219, 42255, 42291, 42328, 42364, 42400, 42437, 
    42473, 42509, 42546, 42582, 42618, 42655, 42691, 42727, 42764, 42800, 
    42837, 42873, 42910, 42946, 42983, 43020, 43056, 43093, 43130, 43167, 
    43204, 43241, 43277, 43314, 43351, 43388, 43425, 43462, 43499, 43536, 
    43573, 43610, 43647, 43684, 43721, 43758, 43794, 43831, 43868, 43905, 
    43942, 43979, 44015, 44052, 44089, 44125, 44162, 44199, 44235, 44272, 
    44308, 44345, 44381, 44418, 44455, 44492, 44528, 44565, 44602, 44639, 
    44676, 44713, 44751, 44788, 44825, 44863, 44900, 44938, 44975, 45012, 
    45050, 45087, 45125, 45162, 45199, 45236, 45273, 45309, 45346, 45382, 
    45418, 45454, 45490, 45526, 45561, 45597, 45632, 45667, 45702, 45737, 
    45772, 45807, 45842, 45877, 45913, 45948, 45983, 46019, 46054, 46090, 
    46126, 46162, 46198, 46234, 46270, 46307, 46344, 46381, 46418, 46455, 
    46492, 46529, 46567, 46604, 46642, 46680, 46717, 46755, 46793, 46830, 
    46868, 46905, 46943, 46980, 47018, 47055, 47092, 47130, 47167, 47203, 
    47240, 47277, 47313, 47350, 47386, 47422, 47458, 47494, 47530, 47566, 
    47601, 47637, 47673, 47708, 47744, 47779, 47815, 47851, 47886, 47922, 
    47958, 47993, 48029, 48065, 48100, 48136, 48172, 48208, 48244, 48280, 
    48316, 48352, 48388, 48424, 48460, 48496, 48532, 48569, 48605, 48641, 
    48678, 48714, 48751, 48787, 48824, 48861, 48898, 48935, 48972, 49009, 
    49046, 49084, 49121, 49159, 49196, 49234, 49271, 49309, 49346, 49383, 
    49421, 49458, 49496, 49533, 49570, 49607, 49644, 49681, 49718, 49755, 
    49792, 49829, 49866, 49903, 49939, 49976, 50013, 50050, 50086, 50123, 
    50160, 50196, 50233, 50270, 50306, 50343, 50379, 50416, 50453, 50489, 
    50525, 50562, 50598, 50634, 50671, 50707, 50743, 50779, 50815, 50851, 
    50887, 50923, 50959, 50994, 51030, 51066, 51102, 51138, 51174, 51210, 
    51246, 51282, 51318, 51354, 51390, 51426, 51462, 51498, 51534, 51570, 
    51606, 51642, 51678, 51714, 51749, 51785, 51821, 51856, 51892, 51927, 
    51963, 51998, 52034, 52069, 52105, 52140, 52176, 52212, 52247, 52283, 
    52319, 52354, 52390, 52426, 52462, 52498, 52534, 52569, 52605, 52641, 
    52677, 52713, 52749, 52786, 52822, 52858, 52894, 52930, 52966, 53003, 
    53039, 53076, 53112, 53149, 53185, 53222, 53259, 53295, 53332, 53369, 
    53405, 53442, 53479, 53515, 53552, 53588, 53625, 53661, 53698, 53734, 
    53770, 53806, 53843, 53879, 53915, 53951, 53987, 54023, 54060, 54096, 
    54132, 54168, 54204, 54240, 54277, 54313, 54349, 54385, 54422, 54458, 
    54494, 54531, 54567, 54603, 54640, 54676, 54712, 54749, 54785, 54821, 
    54858, 54894, 54930, 54967, 55003, 55039, 55076, 55112, 55148, 55185, 
    55221, 55257, 55293, 55330, 55366, 55402, 55438, 55475, 55511, 55547, 
    55583, 55619, 55655, 55691, 55727, 55763, 55799, 55835, 55871, 55907, 
    55943, 55979, 56015, 56051, 56087, 56123, 56159, 56195, 56231, 56268, 
    56304, 56341, 56377, 56414, 56451, 56488, 56524, 56561, 56599, 56636, 
    56673, 56710, 56747, 56784, 56821, 56858, 56895, 56932, 56969, 57006, 
    57043, 57079, 57116, 57152, 57188, 57225, 57261, 57297, 57333, 57369, 
    57405, 57441, 57476, 57512, 57548, 57584, 57620, 57656, 57691, 57727, 
    57763, 57799, 57835, 57871, 57907, 57943, 57979, 58015, 58051, 58087, 
    58122, 58158, 58194, 58230, 58266, 58302, 58338, 58374, 58410, 58446, 
    58482, 58518, 58554, 58590, 58626, 58662, 58699, 58735, 58771, 58807, 
    58843, 58879, 58916, 58952, 58988, 59025, 59061, 59097, 59134, 59170, 
    59207, 59244, 59280, 59317, 59353, 59390, 59427, 59463 ;

 geop_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 press =
  1022.9, 1022.7, 1022.6, 1022.4, 1022.2, 1022, 1021.8, 1021.6, 1021.5, 
    1021.3, 1021.1, 1020.9, 1020.6, 1020.4, 1020.1, 1019.9, 1019.6, 1019.3, 
    1019, 1018.6, 1018.3, 1017.9, 1017.5, 1017.1, 1016.7, 1016.3, 1015.9, 
    1015.5, 1015, 1014.6, 1014.2, 1013.7, 1013.3, 1012.8, 1012.4, 1011.9, 
    1011.4, 1011, 1010.5, 1010, 1009.5, 1009, 1008.5, 1007.9, 1007.4, 1006.9, 
    1006.4, 1005.9, 1005.3, 1004.8, 1004.3, 1003.8, 1003.3, 1002.8, 1002.3, 
    1001.8, 1001.3, 1000.8, 1000.3, 999.81, 999.32, 998.82, 998.32, 997.81, 
    997.31, 996.8, 996.3, 995.79, 995.29, 994.79, 994.29, 993.79, 993.29, 
    992.8, 992.31, 991.83, 991.35, 990.87, 990.39, 989.92, 989.44, 988.97, 
    988.5, 988.04, 987.57, 987.09, 986.62, 986.14, 985.66, 985.18, 984.7, 
    984.22, 983.74, 983.25, 982.76, 982.27, 981.78, 981.28, 980.79, 980.29, 
    979.8, 979.3, 978.8, 978.31, 977.81, 977.31, 976.81, 976.31, 975.81, 
    975.3, 974.8, 974.3, 973.8, 973.3, 972.79, 972.29, 971.79, 971.29, 
    970.78, 970.28, 969.79, 969.29, 968.8, 968.31, 967.82, 967.33, 966.85, 
    966.36, 965.88, 965.4, 964.92, 964.43, 963.95, 963.47, 962.99, 962.51, 
    962.03, 961.55, 961.07, 960.59, 960.1, 959.62, 959.14, 958.66, 958.17, 
    957.69, 957.21, 956.73, 956.25, 955.77, 955.29, 954.81, 954.33, 953.85, 
    953.37, 952.89, 952.4, 951.92, 951.44, 950.95, 950.46, 949.97, 949.47, 
    948.97, 948.47, 947.97, 947.46, 946.95, 946.44, 945.92, 945.41, 944.89, 
    944.36, 943.84, 943.31, 942.79, 942.25, 941.72, 941.19, 940.65, 940.1, 
    939.55, 939, 938.44, 937.88, 937.3, 936.71, 936.12, 935.51, 934.9, 
    934.27, 933.62, 932.97, 932.32, 931.67, 931.01, 930.36, 929.71, 929.07, 
    928.43, 927.79, 927.16, 926.54, 925.91, 925.28, 924.65, 924.03, 923.4, 
    922.77, 922.14, 921.52, 920.89, 920.27, 919.65, 919.03, 918.41, 917.81, 
    917.22, 916.63, 916.04, 915.47, 914.89, 914.33, 913.77, 913.22, 912.69, 
    912.17, 911.66, 911.16, 910.68, 910.21, 909.74, 909.27, 908.81, 908.34, 
    907.87, 907.4, 906.93, 906.45, 905.96, 905.48, 904.99, 904.51, 904.04, 
    903.57, 903.1, 902.63, 902.17, 901.71, 901.26, 900.81, 900.37, 899.93, 
    899.5, 899.06, 898.62, 898.18, 897.74, 897.31, 896.87, 896.44, 896.01, 
    895.6, 895.18, 894.77, 894.36, 893.95, 893.54, 893.14, 892.74, 892.35, 
    891.96, 891.57, 891.18, 890.8, 890.42, 890.05, 889.68, 889.32, 888.96, 
    888.6, 888.24, 887.88, 887.53, 887.18, 886.82, 886.47, 886.12, 885.76, 
    885.4, 885.04, 884.68, 884.31, 883.95, 883.59, 883.23, 882.87, 882.5, 
    882.14, 881.77, 881.39, 881.01, 880.63, 880.24, 879.85, 879.46, 879.06, 
    878.67, 878.27, 877.88, 877.48, 877.09, 876.69, 876.29, 875.9, 875.51, 
    875.11, 874.72, 874.33, 873.94, 873.55, 873.16, 872.77, 872.38, 871.98, 
    871.58, 871.18, 870.78, 870.38, 869.98, 869.59, 869.19, 868.8, 868.42, 
    868.03, 867.65, 867.27, 866.9, 866.53, 866.16, 865.8, 865.45, 865.1, 
    864.75, 864.4, 864.05, 863.69, 863.34, 862.99, 862.63, 862.28, 861.92, 
    861.56, 861.19, 860.83, 860.46, 860.09, 859.72, 859.35, 858.98, 858.61, 
    858.24, 857.87, 857.51, 857.14, 856.78, 856.42, 856.06, 855.69, 855.32, 
    854.95, 854.58, 854.2, 853.82, 853.44, 853.05, 852.67, 852.28, 851.88, 
    851.49, 851.09, 850.69, 850.29, 849.89, 849.49, 849.09, 848.69, 848.29, 
    847.89, 847.49, 847.09, 846.69, 846.29, 845.89, 845.49, 845.08, 844.68, 
    844.27, 843.87, 843.46, 843.06, 842.66, 842.25, 841.85, 841.45, 841.05, 
    840.66, 840.26, 839.86, 839.47, 839.07, 838.68, 838.29, 837.9, 837.51, 
    837.12, 836.72, 836.33, 835.94, 835.55, 835.16, 834.77, 834.38, 833.99, 
    833.6, 833.21, 832.82, 832.43, 832.05, 831.66, 831.28, 830.89, 830.51, 
    830.12, 829.74, 829.36, 828.98, 828.59, 828.21, 827.82, 827.44, 827.05, 
    826.66, 826.27, 825.88, 825.5, 825.11, 824.72, 824.33, 823.95, 823.56, 
    823.17, 822.79, 822.4, 822.02, 821.63, 821.25, 820.87, 820.49, 820.1, 
    819.72, 819.34, 818.96, 818.58, 818.2, 817.81, 817.43, 817.04, 816.66, 
    816.28, 815.9, 815.52, 815.14, 814.76, 814.38, 814, 813.63, 813.26, 
    812.88, 812.51, 812.14, 811.77, 811.4, 811.03, 810.66, 810.28, 809.91, 
    809.53, 809.16, 808.78, 808.4, 808.02, 807.64, 807.25, 806.87, 806.49, 
    806.11, 805.72, 805.34, 804.96, 804.57, 804.19, 803.81, 803.43, 803.05, 
    802.67, 802.29, 801.91, 801.53, 801.15, 800.77, 800.39, 800.01, 799.62, 
    799.24, 798.85, 798.47, 798.08, 797.7, 797.31, 796.93, 796.54, 796.16, 
    795.77, 795.39, 795, 794.62, 794.24, 793.86, 793.48, 793.1, 792.71, 
    792.33, 791.95, 791.57, 791.19, 790.81, 790.43, 790.04, 789.66, 789.28, 
    788.9, 788.52, 788.14, 787.76, 787.38, 787, 786.62, 786.24, 785.86, 
    785.48, 785.1, 784.73, 784.35, 783.97, 783.59, 783.22, 782.84, 782.47, 
    782.09, 781.72, 781.34, 780.97, 780.59, 780.22, 779.85, 779.48, 779.1, 
    778.73, 778.36, 777.99, 777.61, 777.24, 776.87, 776.49, 776.12, 775.74, 
    775.37, 774.99, 774.62, 774.24, 773.86, 773.48, 773.1, 772.72, 772.35, 
    771.97, 771.59, 771.21, 770.83, 770.45, 770.07, 769.69, 769.32, 768.94, 
    768.56, 768.18, 767.8, 767.43, 767.05, 766.67, 766.29, 765.92, 765.54, 
    765.16, 764.78, 764.41, 764.03, 763.65, 763.28, 762.91, 762.53, 762.16, 
    761.79, 761.42, 761.05, 760.69, 760.32, 759.96, 759.59, 759.23, 758.87, 
    758.5, 758.14, 757.78, 757.42, 757.06, 756.7, 756.34, 755.98, 755.61, 
    755.25, 754.89, 754.53, 754.17, 753.8, 753.44, 753.08, 752.71, 752.35, 
    751.99, 751.63, 751.27, 750.91, 750.55, 750.19, 749.84, 749.48, 749.12, 
    748.77, 748.41, 748.06, 747.7, 747.35, 746.99, 746.64, 746.29, 745.94, 
    745.58, 745.23, 744.88, 744.52, 744.17, 743.82, 743.47, 743.11, 742.76, 
    742.41, 742.06, 741.71, 741.36, 741, 740.65, 740.31, 739.96, 739.61, 
    739.27, 738.92, 738.58, 738.23, 737.89, 737.54, 737.2, 736.85, 736.51, 
    736.16, 735.81, 735.46, 735.11, 734.76, 734.41, 734.05, 733.7, 733.34, 
    732.99, 732.63, 732.27, 731.91, 731.55, 731.19, 730.83, 730.47, 730.1, 
    729.74, 729.38, 729.02, 728.66, 728.3, 727.94, 727.58, 727.22, 726.86, 
    726.51, 726.15, 725.79, 725.43, 725.08, 724.72, 724.36, 724.01, 723.65, 
    723.29, 722.94, 722.58, 722.23, 721.87, 721.52, 721.17, 720.82, 720.47, 
    720.11, 719.77, 719.42, 719.07, 718.72, 718.38, 718.03, 717.68, 717.34, 
    716.99, 716.65, 716.31, 715.97, 715.63, 715.29, 714.95, 714.61, 714.27, 
    713.92, 713.58, 713.24, 712.91, 712.57, 712.23, 711.89, 711.55, 711.21, 
    710.87, 710.53, 710.19, 709.86, 709.52, 709.18, 708.85, 708.51, 708.18, 
    707.84, 707.51, 707.17, 706.83, 706.49, 706.15, 705.81, 705.46, 705.11, 
    704.76, 704.4, 704.05, 703.69, 703.34, 702.98, 702.62, 702.26, 701.89, 
    701.53, 701.16, 700.79, 700.43, 700.05, 699.68, 699.31, 698.93, 698.56, 
    698.18, 697.8, 697.42, 697.04, 696.65, 696.27, 695.88, 695.49, 695.1, 
    694.7, 694.31, 693.91, 693.51, 693.12, 692.72, 692.32, 691.92, 691.52, 
    691.12, 690.72, 690.32, 689.92, 689.52, 689.12, 688.72, 688.33, 687.93, 
    687.53, 687.14, 686.74, 686.34, 685.95, 685.56, 685.16, 684.77, 684.38, 
    683.99, 683.6, 683.22, 682.83, 682.45, 682.07, 681.69, 681.31, 680.94, 
    680.56, 680.19, 679.82, 679.46, 679.09, 678.73, 678.38, 678.02, 677.67, 
    677.32, 676.98, 676.63, 676.29, 675.95, 675.62, 675.29, 674.96, 674.63, 
    674.3, 673.97, 673.64, 673.32, 673, 672.67, 672.35, 672.04, 671.72, 
    671.4, 671.09, 670.77, 670.45, 670.14, 669.83, 669.51, 669.2, 668.88, 
    668.57, 668.26, 667.94, 667.63, 667.31, 667, 666.68, 666.37, 666.05, 
    665.74, 665.42, 665.11, 664.79, 664.48, 664.16, 663.84, 663.53, 663.21, 
    662.9, 662.58, 662.27, 661.96, 661.64, 661.33, 661.02, 660.71, 660.39, 
    660.08, 659.77, 659.46, 659.15, 658.84, 658.53, 658.22, 657.91, 657.6, 
    657.29, 656.98, 656.67, 656.36, 656.05, 655.75, 655.44, 655.13, 654.82, 
    654.52, 654.21, 653.91, 653.6, 653.3, 653, 652.7, 652.39, 652.09, 651.79, 
    651.49, 651.19, 650.9, 650.6, 650.3, 650, 649.7, 649.41, 649.11, 648.81, 
    648.51, 648.22, 647.92, 647.62, 647.33, 647.03, 646.74, 646.44, 646.14, 
    645.85, 645.55, 645.26, 644.96, 644.67, 644.38, 644.08, 643.79, 643.5, 
    643.21, 642.91, 642.62, 642.33, 642.03, 641.74, 641.45, 641.15, 640.86, 
    640.56, 640.27, 639.98, 639.68, 639.39, 639.1, 638.81, 638.51, 638.22, 
    637.93, 637.64, 637.35, 637.06, 636.77, 636.48, 636.19, 635.9, 635.61, 
    635.32, 635.03, 634.74, 634.45, 634.16, 633.87, 633.58, 633.29, 633, 
    632.71, 632.42, 632.13, 631.84, 631.55, 631.26, 630.97, 630.68, 630.39, 
    630.1, 629.81, 629.52, 629.22, 628.93, 628.64, 628.35, 628.06, 627.77, 
    627.47, 627.18, 626.89, 626.59, 626.3, 626.01, 625.71, 625.42, 625.13, 
    624.83, 624.54, 624.24, 623.95, 623.65, 623.36, 623.06, 622.77, 622.48, 
    622.18, 621.89, 621.6, 621.3, 621.01, 620.72, 620.43, 620.14, 619.85, 
    619.56, 619.27, 618.97, 618.68, 618.39, 618.1, 617.82, 617.53, 617.24, 
    616.95, 616.66, 616.37, 616.08, 615.79, 615.5, 615.21, 614.93, 614.64, 
    614.35, 614.07, 613.78, 613.5, 613.21, 612.93, 612.65, 612.36, 612.08, 
    611.8, 611.52, 611.23, 610.95, 610.67, 610.39, 610.1, 609.82, 609.54, 
    609.26, 608.97, 608.69, 608.41, 608.13, 607.84, 607.56, 607.28, 607, 
    606.72, 606.44, 606.16, 605.88, 605.6, 605.32, 605.04, 604.76, 604.48, 
    604.2, 603.92, 603.64, 603.36, 603.08, 602.8, 602.51, 602.23, 601.95, 
    601.67, 601.39, 601.11, 600.83, 600.55, 600.27, 599.99, 599.7, 599.42, 
    599.14, 598.86, 598.58, 598.3, 598.01, 597.73, 597.45, 597.17, 596.89, 
    596.6, 596.32, 596.04, 595.76, 595.48, 595.19, 594.91, 594.63, 594.35, 
    594.07, 593.79, 593.51, 593.23, 592.95, 592.67, 592.39, 592.11, 591.83, 
    591.55, 591.27, 590.99, 590.71, 590.43, 590.16, 589.88, 589.6, 589.33, 
    589.05, 588.77, 588.5, 588.22, 587.95, 587.68, 587.4, 587.13, 586.86, 
    586.59, 586.32, 586.04, 585.77, 585.5, 585.23, 584.96, 584.69, 584.42, 
    584.14, 583.87, 583.6, 583.33, 583.07, 582.8, 582.53, 582.26, 581.99, 
    581.72, 581.45, 581.18, 580.91, 580.65, 580.38, 580.11, 579.84, 579.57, 
    579.3, 579.04, 578.77, 578.5, 578.23, 577.96, 577.69, 577.43, 577.16, 
    576.89, 576.62, 576.35, 576.08, 575.81, 575.54, 575.27, 575, 574.73, 
    574.46, 574.19, 573.92, 573.65, 573.38, 573.11, 572.84, 572.58, 572.31, 
    572.04, 571.77, 571.5, 571.23, 570.96, 570.7, 570.43, 570.16, 569.89, 
    569.62, 569.35, 569.09, 568.82, 568.55, 568.28, 568.01, 567.74, 567.48, 
    567.21, 566.94, 566.67, 566.4, 566.14, 565.87, 565.6, 565.34, 565.07, 
    564.8, 564.54, 564.27, 564.01, 563.74, 563.48, 563.21, 562.95, 562.68, 
    562.42, 562.16, 561.89, 561.63, 561.36, 561.1, 560.84, 560.58, 560.31, 
    560.05, 559.79, 559.52, 559.26, 559, 558.74, 558.48, 558.22, 557.96, 
    557.7, 557.44, 557.18, 556.92, 556.66, 556.4, 556.15, 555.89, 555.63, 
    555.37, 555.11, 554.86, 554.6, 554.34, 554.08, 553.82, 553.56, 553.3, 
    553.04, 552.78, 552.52, 552.26, 552.01, 551.75, 551.49, 551.23, 550.97, 
    550.71, 550.45, 550.19, 549.92, 549.66, 549.4, 549.14, 548.88, 548.62, 
    548.36, 548.1, 547.84, 547.58, 547.32, 547.06, 546.8, 546.54, 546.28, 
    546.02, 545.76, 545.5, 545.24, 544.98, 544.72, 544.46, 544.2, 543.94, 
    543.68, 543.42, 543.16, 542.9, 542.65, 542.39, 542.13, 541.87, 541.61, 
    541.35, 541.09, 540.84, 540.58, 540.33, 540.07, 539.81, 539.56, 539.3, 
    539.04, 538.79, 538.53, 538.27, 538.02, 537.76, 537.51, 537.25, 536.99, 
    536.74, 536.48, 536.23, 535.97, 535.72, 535.46, 535.21, 534.95, 534.7, 
    534.45, 534.19, 533.94, 533.69, 533.43, 533.18, 532.93, 532.67, 532.42, 
    532.17, 531.91, 531.66, 531.41, 531.16, 530.9, 530.65, 530.4, 530.15, 
    529.89, 529.64, 529.39, 529.14, 528.88, 528.63, 528.38, 528.13, 527.88, 
    527.63, 527.38, 527.12, 526.87, 526.62, 526.37, 526.12, 525.87, 525.62, 
    525.36, 525.11, 524.86, 524.61, 524.36, 524.11, 523.86, 523.61, 523.36, 
    523.11, 522.85, 522.6, 522.35, 522.1, 521.85, 521.6, 521.35, 521.1, 
    520.85, 520.6, 520.35, 520.1, 519.85, 519.6, 519.36, 519.11, 518.86, 
    518.61, 518.37, 518.12, 517.87, 517.62, 517.38, 517.13, 516.88, 516.64, 
    516.39, 516.15, 515.9, 515.66, 515.41, 515.17, 514.93, 514.68, 514.44, 
    514.2, 513.95, 513.71, 513.47, 513.23, 512.99, 512.74, 512.5, 512.26, 
    512.02, 511.78, 511.54, 511.3, 511.06, 510.82, 510.58, 510.34, 510.1, 
    509.86, 509.62, 509.38, 509.14, 508.9, 508.66, 508.42, 508.18, 507.94, 
    507.7, 507.46, 507.22, 506.98, 506.74, 506.5, 506.26, 506.02, 505.78, 
    505.54, 505.3, 505.07, 504.83, 504.59, 504.35, 504.11, 503.87, 503.63, 
    503.39, 503.15, 502.91, 502.67, 502.43, 502.19, 501.95, 501.72, 501.48, 
    501.24, 501, 500.76, 500.53, 500.29, 500.05, 499.81, 499.58, 499.34, 
    499.1, 498.86, 498.63, 498.39, 498.15, 497.92, 497.68, 497.44, 497.21, 
    496.97, 496.74, 496.5, 496.27, 496.03, 495.8, 495.56, 495.32, 495.09, 
    494.85, 494.62, 494.38, 494.15, 493.91, 493.68, 493.44, 493.21, 492.97, 
    492.74, 492.5, 492.27, 492.03, 491.79, 491.56, 491.32, 491.09, 490.85, 
    490.62, 490.38, 490.15, 489.91, 489.68, 489.44, 489.21, 488.98, 488.74, 
    488.51, 488.27, 488.04, 487.81, 487.57, 487.34, 487.1, 486.87, 486.64, 
    486.41, 486.17, 485.94, 485.71, 485.48, 485.25, 485.02, 484.78, 484.55, 
    484.32, 484.09, 483.86, 483.63, 483.4, 483.17, 482.94, 482.71, 482.48, 
    482.25, 482.02, 481.79, 481.56, 481.33, 481.1, 480.87, 480.64, 480.41, 
    480.18, 479.96, 479.73, 479.5, 479.27, 479.04, 478.81, 478.59, 478.36, 
    478.13, 477.9, 477.67, 477.45, 477.22, 476.99, 476.76, 476.53, 476.31, 
    476.08, 475.85, 475.62, 475.4, 475.17, 474.94, 474.72, 474.49, 474.26, 
    474.04, 473.81, 473.58, 473.36, 473.13, 472.91, 472.68, 472.45, 472.23, 
    472, 471.78, 471.55, 471.33, 471.1, 470.88, 470.65, 470.42, 470.2, 
    469.97, 469.75, 469.52, 469.3, 469.07, 468.85, 468.62, 468.4, 468.17, 
    467.95, 467.72, 467.5, 467.28, 467.05, 466.83, 466.6, 466.38, 466.16, 
    465.93, 465.71, 465.49, 465.26, 465.04, 464.82, 464.59, 464.37, 464.15, 
    463.93, 463.7, 463.48, 463.26, 463.03, 462.81, 462.59, 462.36, 462.14, 
    461.92, 461.69, 461.47, 461.25, 461.02, 460.8, 460.58, 460.35, 460.13, 
    459.91, 459.69, 459.46, 459.24, 459.02, 458.79, 458.57, 458.35, 458.12, 
    457.9, 457.68, 457.46, 457.23, 457.01, 456.79, 456.57, 456.34, 456.12, 
    455.9, 455.68, 455.46, 455.24, 455.01, 454.79, 454.57, 454.35, 454.13, 
    453.91, 453.68, 453.46, 453.24, 453.02, 452.8, 452.58, 452.36, 452.14, 
    451.92, 451.7, 451.48, 451.27, 451.05, 450.83, 450.61, 450.39, 450.17, 
    449.96, 449.74, 449.52, 449.3, 449.08, 448.87, 448.65, 448.43, 448.21, 
    448, 447.78, 447.56, 447.35, 447.13, 446.91, 446.7, 446.48, 446.27, 
    446.05, 445.84, 445.62, 445.41, 445.19, 444.98, 444.77, 444.55, 444.34, 
    444.12, 443.91, 443.7, 443.48, 443.27, 443.05, 442.84, 442.62, 442.41, 
    442.19, 441.98, 441.77, 441.55, 441.34, 441.12, 440.91, 440.7, 440.49, 
    440.27, 440.06, 439.85, 439.63, 439.42, 439.21, 439, 438.78, 438.57, 
    438.36, 438.14, 437.93, 437.72, 437.51, 437.29, 437.08, 436.87, 436.65, 
    436.44, 436.23, 436.02, 435.8, 435.59, 435.38, 435.17, 434.96, 434.74, 
    434.53, 434.32, 434.11, 433.9, 433.69, 433.47, 433.26, 433.05, 432.84, 
    432.63, 432.42, 432.2, 431.99, 431.78, 431.57, 431.36, 431.15, 430.93, 
    430.72, 430.51, 430.3, 430.09, 429.88, 429.67, 429.46, 429.24, 429.03, 
    428.82, 428.61, 428.4, 428.19, 427.98, 427.77, 427.56, 427.35, 427.14, 
    426.93, 426.71, 426.5, 426.3, 426.09, 425.88, 425.67, 425.46, 425.25, 
    425.04, 424.83, 424.62, 424.41, 424.2, 423.99, 423.78, 423.58, 423.37, 
    423.16, 422.95, 422.74, 422.54, 422.33, 422.12, 421.92, 421.71, 421.51, 
    421.3, 421.09, 420.89, 420.68, 420.48, 420.27, 420.07, 419.87, 419.66, 
    419.46, 419.25, 419.05, 418.85, 418.64, 418.44, 418.24, 418.04, 417.83, 
    417.63, 417.43, 417.23, 417.03, 416.82, 416.62, 416.42, 416.22, 416.02, 
    415.82, 415.62, 415.42, 415.22, 415.02, 414.82, 414.62, 414.43, 414.23, 
    414.03, 413.83, 413.63, 413.43, 413.23, 413.03, 412.83, 412.63, 412.43, 
    412.23, 412.03, 411.83, 411.64, 411.44, 411.24, 411.04, 410.84, 410.64, 
    410.44, 410.24, 410.04, 409.84, 409.65, 409.45, 409.25, 409.05, 408.85, 
    408.65, 408.45, 408.25, 408.05, 407.85, 407.65, 407.45, 407.25, 407.05, 
    406.85, 406.66, 406.46, 406.26, 406.06, 405.86, 405.66, 405.46, 405.26, 
    405.06, 404.87, 404.67, 404.47, 404.27, 404.07, 403.87, 403.67, 403.48, 
    403.28, 403.08, 402.88, 402.68, 402.48, 402.28, 402.08, 401.89, 401.69, 
    401.49, 401.29, 401.09, 400.89, 400.7, 400.5, 400.3, 400.1, 399.91, 
    399.71, 399.51, 399.31, 399.11, 398.92, 398.72, 398.52, 398.32, 398.13, 
    397.93, 397.73, 397.53, 397.33, 397.14, 396.94, 396.74, 396.55, 396.35, 
    396.15, 395.96, 395.76, 395.56, 395.37, 395.17, 394.97, 394.78, 394.58, 
    394.39, 394.19, 393.99, 393.8, 393.6, 393.41, 393.21, 393.02, 392.82, 
    392.62, 392.43, 392.23, 392.04, 391.84, 391.65, 391.45, 391.26, 391.06, 
    390.87, 390.67, 390.48, 390.29, 390.09, 389.9, 389.71, 389.52, 389.32, 
    389.13, 388.93, 388.74, 388.55, 388.36, 388.16, 387.97, 387.78, 387.58, 
    387.39, 387.2, 387.01, 386.81, 386.62, 386.43, 386.24, 386.05, 385.85, 
    385.66, 385.47, 385.28, 385.09, 384.9, 384.71, 384.52, 384.33, 384.14, 
    383.95, 383.76, 383.57, 383.38, 383.18, 382.99, 382.8, 382.61, 382.42, 
    382.23, 382.04, 381.85, 381.66, 381.47, 381.28, 381.09, 380.9, 380.71, 
    380.52, 380.33, 380.14, 379.95, 379.76, 379.57, 379.38, 379.19, 379, 
    378.81, 378.63, 378.44, 378.25, 378.06, 377.87, 377.68, 377.5, 377.31, 
    377.12, 376.93, 376.74, 376.55, 376.37, 376.18, 375.99, 375.8, 375.62, 
    375.43, 375.24, 375.05, 374.87, 374.68, 374.5, 374.31, 374.12, 373.94, 
    373.75, 373.57, 373.38, 373.19, 373.01, 372.82, 372.64, 372.45, 372.27, 
    372.08, 371.9, 371.71, 371.53, 371.34, 371.16, 370.97, 370.79, 370.6, 
    370.42, 370.23, 370.05, 369.87, 369.68, 369.5, 369.32, 369.13, 368.95, 
    368.76, 368.58, 368.4, 368.21, 368.03, 367.85, 367.66, 367.48, 367.3, 
    367.11, 366.93, 366.75, 366.56, 366.38, 366.2, 366.02, 365.84, 365.65, 
    365.47, 365.29, 365.11, 364.93, 364.74, 364.56, 364.38, 364.2, 364.02, 
    363.84, 363.66, 363.47, 363.29, 363.11, 362.93, 362.75, 362.56, 362.38, 
    362.2, 362.02, 361.84, 361.66, 361.47, 361.29, 361.11, 360.93, 360.75, 
    360.57, 360.39, 360.21, 360.03, 359.85, 359.67, 359.49, 359.31, 359.13, 
    358.95, 358.77, 358.59, 358.41, 358.23, 358.05, 357.87, 357.69, 357.51, 
    357.33, 357.15, 356.97, 356.79, 356.61, 356.43, 356.25, 356.07, 355.89, 
    355.71, 355.54, 355.36, 355.18, 355, 354.82, 354.65, 354.47, 354.29, 
    354.11, 353.94, 353.76, 353.58, 353.4, 353.23, 353.05, 352.87, 352.7, 
    352.52, 352.34, 352.17, 351.99, 351.81, 351.64, 351.46, 351.28, 351.11, 
    350.93, 350.76, 350.58, 350.4, 350.23, 350.05, 349.88, 349.7, 349.53, 
    349.35, 349.18, 349, 348.83, 348.65, 348.48, 348.31, 348.13, 347.96, 
    347.78, 347.61, 347.43, 347.26, 347.09, 346.91, 346.74, 346.56, 346.39, 
    346.21, 346.04, 345.87, 345.69, 345.52, 345.35, 345.18, 345, 344.83, 
    344.66, 344.48, 344.31, 344.14, 343.97, 343.8, 343.63, 343.45, 343.28, 
    343.11, 342.94, 342.77, 342.59, 342.42, 342.25, 342.08, 341.91, 341.74, 
    341.57, 341.39, 341.22, 341.05, 340.88, 340.71, 340.54, 340.37, 340.2, 
    340.02, 339.85, 339.68, 339.51, 339.34, 339.17, 339, 338.83, 338.66, 
    338.49, 338.31, 338.14, 337.97, 337.8, 337.63, 337.46, 337.29, 337.11, 
    336.94, 336.77, 336.6, 336.43, 336.26, 336.09, 335.92, 335.75, 335.59, 
    335.42, 335.25, 335.08, 334.91, 334.74, 334.57, 334.4, 334.23, 334.06, 
    333.89, 333.73, 333.56, 333.39, 333.22, 333.05, 332.88, 332.72, 332.55, 
    332.38, 332.21, 332.05, 331.88, 331.71, 331.55, 331.38, 331.21, 331.05, 
    330.88, 330.71, 330.55, 330.38, 330.22, 330.05, 329.88, 329.72, 329.55, 
    329.39, 329.22, 329.05, 328.89, 328.72, 328.55, 328.39, 328.22, 328.05, 
    327.89, 327.72, 327.56, 327.39, 327.22, 327.06, 326.89, 326.73, 326.56, 
    326.39, 326.23, 326.06, 325.9, 325.73, 325.56, 325.4, 325.23, 325.07, 
    324.9, 324.74, 324.57, 324.41, 324.24, 324.07, 323.91, 323.74, 323.58, 
    323.41, 323.25, 323.08, 322.92, 322.75, 322.59, 322.42, 322.26, 322.09, 
    321.93, 321.76, 321.6, 321.43, 321.27, 321.1, 320.94, 320.77, 320.61, 
    320.45, 320.28, 320.12, 319.95, 319.79, 319.63, 319.47, 319.3, 319.14, 
    318.98, 318.81, 318.65, 318.49, 318.33, 318.16, 318, 317.84, 317.68, 
    317.51, 317.35, 317.19, 317.03, 316.87, 316.7, 316.54, 316.38, 316.22, 
    316.06, 315.9, 315.73, 315.57, 315.41, 315.25, 315.09, 314.93, 314.77, 
    314.61, 314.45, 314.29, 314.13, 313.97, 313.81, 313.65, 313.49, 313.33, 
    313.17, 313.01, 312.85, 312.69, 312.53, 312.37, 312.21, 312.05, 311.89, 
    311.73, 311.57, 311.41, 311.25, 311.09, 310.93, 310.77, 310.62, 310.46, 
    310.3, 310.14, 309.98, 309.82, 309.66, 309.51, 309.35, 309.19, 309.03, 
    308.87, 308.71, 308.55, 308.4, 308.24, 308.08, 307.92, 307.76, 307.6, 
    307.44, 307.28, 307.13, 306.97, 306.81, 306.65, 306.49, 306.33, 306.18, 
    306.02, 305.86, 305.7, 305.54, 305.39, 305.23, 305.07, 304.91, 304.75, 
    304.6, 304.44, 304.28, 304.12, 303.96, 303.81, 303.65, 303.49, 303.33, 
    303.18, 303.02, 302.86, 302.71, 302.55, 302.39, 302.24, 302.08, 301.92, 
    301.77, 301.61, 301.46, 301.3, 301.14, 300.99, 300.83, 300.68, 300.52, 
    300.36, 300.21, 300.05, 299.9, 299.74, 299.59, 299.43, 299.28, 299.12, 
    298.97, 298.81, 298.66, 298.5, 298.35, 298.2, 298.04, 297.89, 297.74, 
    297.58, 297.43, 297.28, 297.12, 296.97, 296.82, 296.67, 296.51, 296.36, 
    296.21, 296.06, 295.9, 295.75, 295.6, 295.45, 295.29, 295.14, 294.99, 
    294.84, 294.69, 294.54, 294.39, 294.23, 294.08, 293.93, 293.78, 293.63, 
    293.48, 293.33, 293.18, 293.03, 292.88, 292.72, 292.57, 292.42, 292.27, 
    292.12, 291.97, 291.82, 291.67, 291.52, 291.37, 291.22, 291.07, 290.92, 
    290.77, 290.62, 290.47, 290.32, 290.17, 290.02, 289.87, 289.72, 289.57, 
    289.42, 289.28, 289.13, 288.98, 288.83, 288.68, 288.53, 288.38, 288.23, 
    288.08, 287.93, 287.79, 287.64, 287.49, 287.34, 287.19, 287.04, 286.9, 
    286.75, 286.6, 286.45, 286.3, 286.15, 286.01, 285.86, 285.71, 285.56, 
    285.41, 285.26, 285.12, 284.97, 284.82, 284.67, 284.52, 284.38, 284.23, 
    284.08, 283.93, 283.78, 283.64, 283.49, 283.34, 283.19, 283.05, 282.9, 
    282.75, 282.6, 282.46, 282.31, 282.16, 282.01, 281.87, 281.72, 281.57, 
    281.43, 281.28, 281.13, 280.99, 280.84, 280.69, 280.55, 280.4, 280.25, 
    280.11, 279.96, 279.81, 279.67, 279.52, 279.37, 279.23, 279.08, 278.93, 
    278.79, 278.64, 278.5, 278.35, 278.2, 278.06, 277.91, 277.76, 277.62, 
    277.47, 277.33, 277.18, 277.03, 276.89, 276.74, 276.6, 276.45, 276.31, 
    276.16, 276.02, 275.87, 275.73, 275.58, 275.44, 275.29, 275.15, 275, 
    274.86, 274.72, 274.57, 274.43, 274.28, 274.14, 274, 273.85, 273.71, 
    273.56, 273.42, 273.28, 273.13, 272.99, 272.85, 272.7, 272.56, 272.42, 
    272.27, 272.13, 271.99, 271.84, 271.7, 271.56, 271.42, 271.27, 271.13, 
    270.99, 270.84, 270.7, 270.56, 270.42, 270.27, 270.13, 269.99, 269.85, 
    269.7, 269.56, 269.42, 269.28, 269.13, 268.99, 268.85, 268.71, 268.57, 
    268.42, 268.28, 268.14, 268, 267.86, 267.72, 267.57, 267.43, 267.29, 
    267.15, 267.01, 266.87, 266.73, 266.59, 266.44, 266.3, 266.16, 266.02, 
    265.88, 265.74, 265.6, 265.46, 265.32, 265.18, 265.04, 264.9, 264.76, 
    264.62, 264.48, 264.34, 264.2, 264.05, 263.91, 263.77, 263.63, 263.49, 
    263.35, 263.21, 263.07, 262.93, 262.8, 262.66, 262.52, 262.38, 262.24, 
    262.1, 261.96, 261.82, 261.68, 261.55, 261.41, 261.27, 261.13, 260.99, 
    260.86, 260.72, 260.58, 260.44, 260.3, 260.17, 260.03, 259.89, 259.75, 
    259.62, 259.48, 259.34, 259.2, 259.07, 258.93, 258.79, 258.65, 258.52, 
    258.38, 258.24, 258.11, 257.97, 257.84, 257.7, 257.56, 257.43, 257.29, 
    257.15, 257.02, 256.88, 256.75, 256.61, 256.47, 256.34, 256.2, 256.07, 
    255.93, 255.79, 255.66, 255.52, 255.39, 255.25, 255.12, 254.98, 254.85, 
    254.71, 254.58, 254.44, 254.31, 254.17, 254.04, 253.91, 253.77, 253.64, 
    253.5, 253.37, 253.23, 253.1, 252.96, 252.83, 252.7, 252.56, 252.43, 
    252.29, 252.16, 252.03, 251.89, 251.76, 251.62, 251.49, 251.36, 251.22, 
    251.09, 250.96, 250.82, 250.69, 250.55, 250.42, 250.29, 250.15, 250.02, 
    249.89, 249.75, 249.62, 249.49, 249.36, 249.22, 249.09, 248.96, 248.83, 
    248.69, 248.56, 248.43, 248.3, 248.16, 248.03, 247.9, 247.77, 247.63, 
    247.5, 247.37, 247.23, 247.1, 246.97, 246.84, 246.71, 246.57, 246.44, 
    246.31, 246.18, 246.05, 245.92, 245.79, 245.65, 245.52, 245.39, 245.26, 
    245.13, 245, 244.87, 244.74, 244.61, 244.48, 244.34, 244.21, 244.08, 
    243.95, 243.82, 243.69, 243.56, 243.43, 243.3, 243.17, 243.04, 242.91, 
    242.78, 242.65, 242.52, 242.39, 242.26, 242.13, 242, 241.87, 241.75, 
    241.62, 241.49, 241.36, 241.23, 241.1, 240.97, 240.84, 240.71, 240.58, 
    240.45, 240.32, 240.19, 240.06, 239.93, 239.81, 239.68, 239.55, 239.42, 
    239.29, 239.16, 239.03, 238.91, 238.78, 238.65, 238.52, 238.39, 238.26, 
    238.14, 238.01, 237.88, 237.75, 237.62, 237.5, 237.37, 237.24, 237.11, 
    236.99, 236.86, 236.73, 236.61, 236.48, 236.35, 236.23, 236.1, 235.97, 
    235.85, 235.72, 235.59, 235.47, 235.34, 235.22, 235.09, 234.96, 234.84, 
    234.71, 234.59, 234.46, 234.34, 234.21, 234.08, 233.96, 233.83, 233.71, 
    233.58, 233.46, 233.33, 233.21, 233.08, 232.96, 232.83, 232.7, 232.58, 
    232.45, 232.33, 232.2, 232.08, 231.95, 231.83, 231.7, 231.57, 231.45, 
    231.32, 231.2, 231.07, 230.95, 230.82, 230.7, 230.57, 230.45, 230.32, 
    230.2, 230.07, 229.95, 229.82, 229.7, 229.57, 229.45, 229.32, 229.2, 
    229.07, 228.95, 228.82, 228.7, 228.57, 228.45, 228.32, 228.2, 228.07, 
    227.95, 227.82, 227.7, 227.57, 227.45, 227.32, 227.2, 227.07, 226.95, 
    226.82, 226.7, 226.58, 226.45, 226.33, 226.2, 226.08, 225.95, 225.83, 
    225.7, 225.58, 225.46, 225.33, 225.21, 225.08, 224.96, 224.84, 224.71, 
    224.59, 224.46, 224.34, 224.22, 224.09, 223.97, 223.85, 223.72, 223.6, 
    223.48, 223.35, 223.23, 223.11, 222.98, 222.86, 222.74, 222.62, 222.49, 
    222.37, 222.25, 222.12, 222, 221.88, 221.75, 221.63, 221.51, 221.39, 
    221.27, 221.14, 221.02, 220.9, 220.78, 220.66, 220.54, 220.41, 220.29, 
    220.17, 220.05, 219.93, 219.81, 219.68, 219.56, 219.44, 219.32, 219.2, 
    219.08, 218.95, 218.83, 218.71, 218.59, 218.47, 218.35, 218.23, 218.11, 
    217.99, 217.86, 217.74, 217.62, 217.5, 217.38, 217.26, 217.14, 217.02, 
    216.9, 216.78, 216.66, 216.54, 216.42, 216.3, 216.18, 216.05, 215.93, 
    215.81, 215.69, 215.57, 215.45, 215.33, 215.21, 215.09, 214.98, 214.86, 
    214.74, 214.62, 214.5, 214.38, 214.26, 214.14, 214.02, 213.9, 213.78, 
    213.66, 213.54, 213.43, 213.31, 213.19, 213.07, 212.95, 212.83, 212.72, 
    212.6, 212.48, 212.36, 212.24, 212.12, 212, 211.89, 211.77, 211.65, 
    211.53, 211.41, 211.3, 211.18, 211.06, 210.94, 210.82, 210.71, 210.59, 
    210.47, 210.36, 210.24, 210.12, 210.01, 209.89, 209.78, 209.66, 209.54, 
    209.43, 209.31, 209.2, 209.08, 208.97, 208.85, 208.74, 208.63, 208.51, 
    208.4, 208.28, 208.17, 208.06, 207.95, 207.83, 207.72, 207.61, 207.5, 
    207.39, 207.27, 207.16, 207.05, 206.94, 206.83, 206.72, 206.61, 206.49, 
    206.38, 206.27, 206.16, 206.05, 205.94, 205.83, 205.72, 205.61, 205.5, 
    205.39, 205.28, 205.17, 205.06, 204.95, 204.84, 204.72, 204.61, 204.5, 
    204.39, 204.28, 204.17, 204.06, 203.95, 203.84, 203.73, 203.62, 203.51, 
    203.4, 203.29, 203.18, 203.07, 202.96, 202.85, 202.74, 202.63, 202.52, 
    202.41, 202.31, 202.2, 202.09, 201.98, 201.87, 201.76, 201.65, 201.54, 
    201.43, 201.33, 201.22, 201.11, 201, 200.89, 200.78, 200.67, 200.57, 
    200.46, 200.35, 200.24, 200.14, 200.03, 199.92, 199.81, 199.7, 199.6, 
    199.49, 199.38, 199.27, 199.17, 199.06, 198.95, 198.84, 198.73, 198.63, 
    198.52, 198.41, 198.3, 198.19, 198.09, 197.98, 197.87, 197.76, 197.65, 
    197.54, 197.43, 197.33, 197.22, 197.11, 197, 196.89, 196.78, 196.67, 
    196.57, 196.46, 196.35, 196.24, 196.13, 196.02, 195.92, 195.81, 195.7, 
    195.59, 195.48, 195.38, 195.27, 195.16, 195.05, 194.95, 194.84, 194.73, 
    194.62, 194.52, 194.41, 194.3, 194.19, 194.09, 193.98, 193.87, 193.77, 
    193.66, 193.56, 193.45, 193.34, 193.24, 193.13, 193.03, 192.92, 192.81, 
    192.71, 192.6, 192.5, 192.39, 192.29, 192.18, 192.08, 191.97, 191.86, 
    191.76, 191.65, 191.55, 191.44, 191.34, 191.23, 191.12, 191.02, 190.91, 
    190.81, 190.7, 190.6, 190.49, 190.39, 190.28, 190.18, 190.07, 189.97, 
    189.86, 189.76, 189.65, 189.55, 189.45, 189.34, 189.24, 189.13, 189.03, 
    188.93, 188.82, 188.72, 188.62, 188.51, 188.41, 188.31, 188.2, 188.1, 
    188, 187.9, 187.79, 187.69, 187.59, 187.49, 187.38, 187.28, 187.18, 
    187.08, 186.98, 186.88, 186.78, 186.68, 186.57, 186.47, 186.37, 186.27, 
    186.17, 186.07, 185.96, 185.86, 185.76, 185.66, 185.56, 185.45, 185.35, 
    185.25, 185.15, 185.05, 184.95, 184.84, 184.74, 184.64, 184.54, 184.44, 
    184.34, 184.24, 184.14, 184.03, 183.93, 183.83, 183.73, 183.63, 183.53, 
    183.43, 183.33, 183.23, 183.13, 183.03, 182.93, 182.83, 182.73, 182.63, 
    182.53, 182.43, 182.33, 182.23, 182.13, 182.03, 181.93, 181.83, 181.73, 
    181.63, 181.53, 181.44, 181.34, 181.24, 181.14, 181.04, 180.94, 180.84, 
    180.74, 180.65, 180.55, 180.45, 180.35, 180.25, 180.15, 180.05, 179.96, 
    179.86, 179.76, 179.66, 179.56, 179.46, 179.37, 179.27, 179.17, 179.07, 
    178.97, 178.88, 178.78, 178.68, 178.58, 178.49, 178.39, 178.29, 178.2, 
    178.1, 178, 177.91, 177.81, 177.72, 177.62, 177.52, 177.43, 177.33, 
    177.24, 177.14, 177.04, 176.95, 176.85, 176.76, 176.66, 176.57, 176.47, 
    176.38, 176.28, 176.18, 176.09, 175.99, 175.9, 175.8, 175.71, 175.61, 
    175.52, 175.43, 175.33, 175.24, 175.14, 175.05, 174.95, 174.86, 174.76, 
    174.67, 174.58, 174.48, 174.39, 174.3, 174.2, 174.11, 174.02, 173.92, 
    173.83, 173.74, 173.64, 173.55, 173.46, 173.37, 173.27, 173.18, 173.09, 
    173, 172.9, 172.81, 172.72, 172.63, 172.54, 172.45, 172.35, 172.26, 
    172.17, 172.08, 171.99, 171.9, 171.81, 171.72, 171.63, 171.53, 171.44, 
    171.35, 171.26, 171.17, 171.08, 170.99, 170.9, 170.8, 170.71, 170.62, 
    170.53, 170.44, 170.35, 170.26, 170.16, 170.07, 169.98, 169.89, 169.8, 
    169.71, 169.62, 169.53, 169.44, 169.35, 169.25, 169.16, 169.07, 168.98, 
    168.89, 168.8, 168.71, 168.62, 168.53, 168.44, 168.35, 168.26, 168.17, 
    168.08, 167.99, 167.9, 167.81, 167.72, 167.63, 167.54, 167.45, 167.36, 
    167.27, 167.18, 167.09, 167, 166.91, 166.82, 166.73, 166.64, 166.55, 
    166.46, 166.37, 166.29, 166.2, 166.11, 166.02, 165.93, 165.84, 165.75, 
    165.66, 165.57, 165.48, 165.4, 165.31, 165.22, 165.13, 165.04, 164.95, 
    164.86, 164.78, 164.69, 164.6, 164.51, 164.42, 164.34, 164.25, 164.16, 
    164.07, 163.99, 163.9, 163.81, 163.72, 163.64, 163.55, 163.46, 163.38, 
    163.29, 163.2, 163.12, 163.03, 162.94, 162.86, 162.77, 162.69, 162.6, 
    162.51, 162.43, 162.34, 162.26, 162.17, 162.08, 162, 161.91, 161.83, 
    161.74, 161.66, 161.57, 161.49, 161.4, 161.31, 161.23, 161.14, 161.06, 
    160.97, 160.89, 160.8, 160.72, 160.63, 160.55, 160.46, 160.38, 160.29, 
    160.21, 160.12, 160.04, 159.95, 159.87, 159.78, 159.7, 159.61, 159.53, 
    159.45, 159.36, 159.28, 159.19, 159.11, 159.02, 158.94, 158.85, 158.77, 
    158.69, 158.6, 158.52, 158.43, 158.35, 158.27, 158.18, 158.1, 158.01, 
    157.93, 157.85, 157.76, 157.68, 157.6, 157.51, 157.43, 157.34, 157.26, 
    157.18, 157.09, 157.01, 156.93, 156.85, 156.76, 156.68, 156.6, 156.51, 
    156.43, 156.35, 156.27, 156.18, 156.1, 156.02, 155.94, 155.85, 155.77, 
    155.69, 155.61, 155.53, 155.44, 155.36, 155.28, 155.2, 155.12, 155.04, 
    154.96, 154.87, 154.79, 154.71, 154.63, 154.55, 154.47, 154.39, 154.31, 
    154.23, 154.15, 154.06, 153.98, 153.9, 153.82, 153.74, 153.66, 153.58, 
    153.5, 153.42, 153.34, 153.26, 153.18, 153.1, 153.02, 152.94, 152.86, 
    152.59, 152.33, 152.07, 151.81, 151.57, 151.32, 151.08, 150.84, 150.61, 
    150.37, 150.13, 149.9, 149.66, 149.41, 149.16, 148.91, 148.65, 148.38, 
    148.11, 147.84, 147.55, 147.26, 146.96, 146.66, 146.36, 146.05, 145.74, 
    145.42, 145.11, 144.79, 144.48, 144.16, 143.85, 143.55, 143.24, 142.94, 
    142.65, 142.35, 142.07, 141.78, 141.5, 141.23, 140.96, 140.69, 140.42, 
    140.15, 139.89, 139.62, 139.36, 139.1, 138.83, 138.56, 138.3, 138.03, 
    137.76, 137.48, 137.21, 136.93, 136.65, 136.37, 136.09, 135.81, 135.52, 
    135.24, 134.95, 134.67, 134.39, 134.1, 133.82, 133.54, 133.26, 132.99, 
    132.71, 132.44, 132.17, 131.9, 131.63, 131.37, 131.1, 130.84, 130.58, 
    130.31, 130.05, 129.79, 129.53, 129.26, 129, 128.73, 128.46, 128.19, 
    127.92, 127.65, 127.38, 127.1, 126.83, 126.55, 126.28, 126, 125.72, 
    125.44, 125.16, 124.88, 124.6, 124.33, 124.05, 123.77, 123.49, 123.22, 
    122.94, 122.66, 122.39, 122.11, 121.84, 121.57, 121.3, 121.03, 120.76, 
    120.49, 120.22, 119.95, 119.69, 119.43, 119.16, 118.9, 118.64, 118.38, 
    118.13, 117.87, 117.62, 117.36, 117.11, 116.86, 116.61, 116.36, 116.11, 
    115.86, 115.61, 115.36, 115.11, 114.86, 114.61, 114.36, 114.11, 113.86, 
    113.6, 113.35, 113.09, 112.83, 112.57, 112.31, 112.05, 111.78, 111.51, 
    111.24, 110.97, 110.69, 110.42, 110.14, 109.86, 109.58, 109.3, 109.02, 
    108.74, 108.46, 108.18, 107.9, 107.62, 107.33, 107.05, 106.77, 106.49, 
    106.22, 105.94, 105.66, 105.38, 105.11, 104.84, 104.56, 104.29, 104.02, 
    103.75, 103.48, 103.21, 102.94, 102.67, 102.41, 102.14, 101.88, 101.61, 
    101.35, 101.08, 100.82, 100.56, 100.3, 100.04, 99.775, 99.515, 99.255, 
    98.995, 98.734, 98.474, 98.213, 97.951, 97.687, 97.423, 97.156, 96.887, 
    96.616, 96.342, 96.065, 95.785, 95.501, 95.214, 94.924, 94.63, 94.332, 
    94.032, 93.728, 93.422, 93.113, 92.802, 92.489, 92.175, 91.859, 91.543, 
    91.226, 90.909, 90.593, 90.277, 89.962, 89.648, 89.335, 89.024, 88.714, 
    88.405, 88.098, 87.793, 87.489, 87.187, 86.887, 86.588, 86.29, 85.994, 
    85.7, 85.407, 85.116, 84.827, 84.54, 84.255, 83.972, 83.692, 83.415, 
    83.14, 82.869, 82.602, 82.337, 82.077, 81.821, 81.568, 81.32, 81.076, 
    80.836, 80.601, 80.369, 80.142, 79.919, 79.699, 79.483, 79.27, 79.06, 
    78.853, 78.649, 78.446, 78.245, 78.046, 77.848, 77.65, 77.453, 77.257, 
    77.06, 76.864, 76.667, 76.47, 76.273, 76.076, 75.878, 75.681, 75.483, 
    75.286, 75.088, 74.891, 74.694, 74.497, 74.3, 74.104, 73.908, 73.711, 
    73.515, 73.318, 73.121, 72.922, 72.723, 72.523, 72.321, 72.118, 71.913, 
    71.706, 71.496, 71.285, 71.071, 70.856, 70.637, 70.417, 70.194, 69.969, 
    69.742, 69.513, 69.281, 69.048, 68.813, 68.576, 68.338, 68.097, 67.856, 
    67.612, 67.368, 67.122, 66.876, 66.628, 66.379, 66.13, 65.881, 65.63, 
    65.38, 65.13, 64.879, 64.629, 64.379, 64.13, 63.881, 63.634, 63.387, 
    63.141, 62.896, 62.653, 62.411, 62.171, 61.933, 61.696, 61.46, 61.227, 
    60.996, 60.766, 60.539, 60.313, 60.09, 59.868, 59.648, 59.431, 59.215, 
    59.001, 58.79, 58.58, 58.372, 58.166, 57.961, 57.759, 57.558, 57.359, 
    57.162, 56.966, 56.771, 56.578, 56.387, 56.196, 56.007, 55.819, 55.632, 
    55.446, 55.262, 55.078, 54.895, 54.713, 54.531, 54.351, 54.171, 53.992, 
    53.814, 53.637, 53.46, 53.284, 53.109, 52.935, 52.761, 52.588, 52.415, 
    52.243, 52.071, 51.899, 51.727, 51.555, 51.382, 51.209, 51.036, 50.862, 
    50.687, 50.511, 50.335, 50.157, 49.978, 49.799, 49.619, 49.437, 49.256, 
    49.073, 48.89, 48.707, 48.524, 48.341, 48.159, 47.976, 47.795, 47.614, 
    47.434, 47.255, 47.077, 46.9, 46.725, 46.551, 46.377, 46.205, 46.035, 
    45.865, 45.696, 45.528, 45.361, 45.194, 45.028, 44.862, 44.697, 44.532, 
    44.368, 44.203, 44.039, 43.875, 43.711, 43.547, 43.383, 43.22, 43.057, 
    42.894, 42.731, 42.568, 42.406, 42.244, 42.082, 41.92, 41.759, 41.597, 
    41.435, 41.273, 41.111, 40.948, 40.785, 40.621, 40.457, 40.292, 40.126, 
    39.959, 39.792, 39.624, 39.455, 39.285, 39.115, 38.945, 38.774, 38.603, 
    38.432, 38.261, 38.091, 37.921, 37.751, 37.582, 37.414, 37.247, 37.081, 
    36.917, 36.754, 36.592, 36.432, 36.273, 36.117, 35.962, 35.809, 35.658, 
    35.509, 35.362, 35.216, 35.073, 34.932, 34.792, 34.654, 34.518, 34.384, 
    34.251, 34.119, 33.989, 33.86, 33.731, 33.604, 33.477, 33.35, 33.223, 
    33.096, 32.969, 32.842, 32.714, 32.586, 32.456, 32.326, 32.195, 32.062, 
    31.929, 31.794, 31.659, 31.522, 31.384, 31.246, 31.106, 30.966, 30.825, 
    30.683, 30.542, 30.399, 30.257, 30.115, 29.972, 29.83, 29.689, 29.548, 
    29.407, 29.267, 29.128, 28.989, 28.851, 28.715, 28.579, 28.444, 28.309, 
    28.176, 28.044, 27.912, 27.781, 27.651, 27.521, 27.392, 27.264, 27.136, 
    27.01, 26.883, 26.758, 26.633, 26.51, 26.387, 26.265, 26.144, 26.024, 
    25.905, 25.788, 25.671, 25.556, 25.443, 25.33, 25.219, 25.109, 25, 
    24.892, 24.786, 24.68, 24.575, 24.471, 24.368, 24.265, 24.163, 24.061, 
    23.959, 23.857, 23.756, 23.654, 23.553, 23.451, 23.349, 23.247, 23.145, 
    23.042, 22.939, 22.836, 22.732, 22.628, 22.524, 22.419, 22.314, 22.209, 
    22.103, 21.997, 21.89, 21.784, 21.676, 21.569, 21.461, 21.354, 21.246, 
    21.138, 21.03, 20.922, 20.815, 20.708, 20.601, 20.494, 20.388, 20.282, 
    20.177, 20.073, 19.969, 19.866, 19.764, 19.662, 19.561, 19.46, 19.361, 
    19.261, 19.163, 19.065, 18.968, 18.871, 18.775, 18.68, 18.586, 18.492, 
    18.398, 18.306, 18.214, 18.122, 18.032, 17.942, 17.852, 17.764, 17.675, 
    17.588, 17.501, 17.414, 17.328, 17.242, 17.157, 17.072, 16.988, 16.904, 
    16.82, 16.737, 16.655, 16.573, 16.491, 16.411, 16.331, 16.251, 16.173, 
    16.095, 16.018, 15.941, 15.865, 15.79, 15.716, 15.642, 15.568, 15.495, 
    15.422, 15.35, 15.278, 15.206, 15.134, 15.062, 14.99, 14.918, 14.846, 
    14.774, 14.702, 14.629, 14.557, 14.484, 14.411, 14.337, 14.264, 14.19, 
    14.116, 14.042, 13.967, 13.893, 13.818, 13.743, 13.668, 13.593, 13.518, 
    13.443, 13.368, 13.294, 13.219, 13.145, 13.071, 12.997, 12.924, 12.851, 
    12.778, 12.706, 12.635, 12.564, 12.494, 12.425, 12.356, 12.287, 12.22, 
    12.153, 12.086, 12.02, 11.955, 11.89, 11.826, 11.762, 11.699, 11.636, 
    11.574, 11.512, 11.451, 11.39, 11.329, 11.269, 11.21, 11.15, 11.091, 
    11.033, 10.975, 10.917, 10.859, 10.802, 10.745, 10.689, 10.632, 10.577, 
    10.521, 10.466, 10.411, 10.356, 10.302, 10.248, 10.194, 10.141, 10.088, 
    10.035, 9.9828, 9.9308, 9.8792, 9.8279, 9.7769, 9.7263, 9.6761, 9.6262, 
    9.5767, 9.5276, 9.4788, 9.4303, 9.3823, 9.3345, 9.2872, 9.2402, 9.1935, 
    9.1472, 9.1012, 9.0555, 9.01, 8.9649, 8.9199, 8.8752, 8.8307, 8.7863, 
    8.742, 8.6979, 8.6538, 8.6098, 8.5659, 8.522, 8.4781, 8.4342, 8.3903, 
    8.3465, 8.3026, 8.2588, 8.2149, 8.1711, 8.1274, 8.0837, 8.0401, 7.9966, 
    7.9532, 7.91, 7.8669, 7.824, 7.7813, 7.7388, 7.6965, 7.6545, 7.6127, 
    7.5712, 7.53, 7.489, 7.4483, 7.4079, 7.3678, 7.3279, 7.2884, 7.2491, 
    7.2101, 7.1713, 7.1328, 7.0946, 7.0567, 7.019, 6.9815, 6.9443, 6.9072, 
    6.8704, 6.8338, 6.7974, 6.7612, 6.7251, 6.6892, 6.6535, 6.6179, 6.5824, 
    6.5471, 6.5118, 6.4768, 6.4418, 6.4069, 6.3722, 6.3377, 6.3032, 6.2689, 
    6.2348, 6.2008, 6.1669, 6.1333, 6.0998, 6.0665, 6.0335, 6.0006, 5.9679, 
    5.9354, 5.9031, 5.871, 5.8391, 5.8074, 5.7759, 5.7446, 5.7135, 5.6825, 
    5.6517, 5.6211, 5.5906, 5.5602, 5.5301, 5.5, 5.4701, 5.4403, 5.4107, 
    5.3812, 5.3518, 5.3226, 5.2935, 5.2646, 5.2358, 5.2071, 5.1786, 5.1503, 
    5.1221, 5.0941, 5.0662, 5.0385, 5.011, 4.9837, 4.9566, 4.9296, 4.9029, 
    4.8763, 4.85, 4.8238, 4.7979, 4.7721, 4.7465, 4.7212, 4.696, 4.671, 
    4.6462, 4.6215, 4.5971, 4.5728, 4.5486, 4.5247, 4.5009, 4.4772, 4.4537, 
    4.4303, 4.4071, 4.3841, 4.3611, 4.3383, 4.3157, 4.2931, 4.2707, 4.2485, 
    4.2263, 4.2043, 4.1824, 4.1606, 4.1389, 4.1173, 4.0959, 4.0745, 4.0532, 
    4.032, 4.0109, 3.9898, 3.9689, 3.948, 3.9272, 3.9065, 3.8859, 3.8653, 
    3.8449, 3.8245, 3.8043, 3.7842, 3.7642, 3.7443, 3.7245, 3.7049, 3.6855, 
    3.6661, 3.647, 3.6279, 3.609, 3.5903, 3.5717, 3.5532, 3.5349, 3.5166, 
    3.4985, 3.4805, 3.4626, 3.4447, 3.427, 3.4093, 3.3917, 3.3741, 3.3567, 
    3.3392, 3.3219, 3.3046, 3.2873, 3.2701, 3.253, 3.236, 3.219, 3.2021, 
    3.1853, 3.1686, 3.1519, 3.1354, 3.1189, 3.1026, 3.0864, 3.0702, 3.0542, 
    3.0383, 3.0225, 3.0069, 2.9913, 2.9759, 2.9606, 2.9454, 2.9304, 2.9155, 
    2.9007, 2.886, 2.8714, 2.857, 2.8427, 2.8284, 2.8143, 2.8003, 2.7865, 
    2.7727, 2.759, 2.7454, 2.7318, 2.7184, 2.705, 2.6917, 2.6785, 2.6653, 
    2.6522, 2.6391, 2.6261, 2.6132, 2.6003, 2.5874, 2.5745, 2.5618, 2.549, 
    2.5363, 2.5236, 2.5109, 2.4983, 2.4857, 2.4731, 2.4606, 2.4481, 2.4356, 
    2.4232, 2.4109, 2.3986, 2.3863, 2.3741, 2.3619, 2.3498, 2.3378, 2.3258, 
    2.3139, 2.3021, 2.2903, 2.2786, 2.267, 2.2555, 2.2441, 2.2327, 2.2214, 
    2.2102, 2.1991, 2.188, 2.177, 2.1662, 2.1553, 2.1446, 2.1339, 2.1233, 
    2.1128, 2.1024, 2.092, 2.0817, 2.0714, 2.0612, 2.0511, 2.0411, 2.0311, 
    2.0212, 2.0113, 2.0015, 1.9918, 1.9822, 1.9726, 1.963, 1.9535, 1.9441, 
    1.9348, 1.9254, 1.9162, 1.907, 1.8978, 1.8887, 1.8796, 1.8706, 1.8616, 
    1.8527, 1.8438, 1.835, 1.8262, 1.8175, 1.8088, 1.8001, 1.7915, 1.783, 
    1.7745, 1.766, 1.7576, 1.7492, 1.7408, 1.7326, 1.7243, 1.7161, 1.708, 
    1.6998, 1.6918, 1.6837, 1.6757, 1.6678, 1.6598, 1.652, 1.6441, 1.6363, 
    1.6285, 1.6208, 1.6131, 1.6055, 1.5979, 1.5903, 1.5828, 1.5753, 1.5678, 
    1.5604, 1.553, 1.5457, 1.5384, 1.5312, 1.524, 1.5168, 1.5097, 1.5026, 
    1.4956, 1.4886, 1.4817, 1.4747, 1.4679, 1.461, 1.4542, 1.4475, 1.4407, 
    1.4341, 1.4274, 1.4208, 1.4143, 1.4077, 1.4012, 1.3948, 1.3884, 1.382, 
    1.3756, 1.3693, 1.363, 1.3567, 1.3505, 1.3443, 1.3381, 1.332, 1.3259, 
    1.3198, 1.3137, 1.3076, 1.3016, 1.2956, 1.2897, 1.2837, 1.2778, 1.2719, 
    1.266, 1.2602, 1.2544, 1.2486, 1.2429, 1.2372, 1.2315, 1.2258, 1.2202, 
    1.2146, 1.209, 1.2035, 1.1979, 1.1925, 1.187, 1.1816, 1.1762, 1.1708, 
    1.1655, 1.1602, 1.155, 1.1497, 1.1445, 1.1393, 1.1342, 1.1291, 1.124, 
    1.119, 1.1139, 1.1089, 1.104, 1.099, 1.0941, 1.0892, 1.0843, 1.0794, 
    1.0746, 1.0697, 1.0649, 1.0601, 1.0553, 1.0505, 1.0457, 1.0409, 1.0362, 
    1.0315, 1.0268, 1.0221, 1.0175, 1.0128, 1.0082, 1.0037, 0.99916, 0.99468, 
    0.99023, 0.98582, 0.98146, 0.97713, 0.97285, 0.9686, 0.9644, 0.96024, 
    0.95612, 0.95203, 0.94798, 0.94396, 0.93998, 0.93602, 0.93208, 0.92817, 
    0.92428, 0.9204, 0.91654, 0.91269, 0.90885, 0.90502, 0.9012, 0.89738, 
    0.89356, 0.88975, 0.88594, 0.88213, 0.87832, 0.87451, 0.8707, 0.8669, 
    0.8631, 0.85931, 0.85552, 0.85173, 0.84796, 0.84419, 0.84043, 0.83669, 
    0.83296, 0.82924, 0.82554, 0.82186, 0.81819, 0.81455, 0.81092, 0.80732, 
    0.80374, 0.80019, 0.79666, 0.79316, 0.78968, 0.78623, 0.78281, 0.77942, 
    0.77605, 0.77271, 0.7694, 0.76611, 0.76285, 0.75962, 0.7564, 0.75322, 
    0.75005, 0.7469, 0.74377, 0.74066, 0.73757, 0.73449, 0.73142, 0.72837, 
    0.72533, 0.7223, 0.71928, 0.71628, 0.71328, 0.7103, 0.70732, 0.70436, 
    0.70141, 0.69846, 0.69553, 0.6926, 0.68969, 0.68679, 0.68389, 0.68101, 
    0.67814, 0.67527, 0.67241, 0.66957, 0.66673, 0.66389, 0.66107, 0.65825, 
    0.65544, 0.65263, 0.64983, 0.64703, 0.64423, 0.64144, 0.63866, 0.63588, 
    0.6331, 0.63033, 0.62756, 0.6248, 0.62205, 0.61931, 0.61658, 0.61385, 
    0.61114, 0.60844, 0.60575, 0.60307, 0.60041, 0.59776, 0.59513, 0.5925, 
    0.5899, 0.58731, 0.58473, 0.58217, 0.57961, 0.57708, 0.57455, 0.57204, 
    0.56954, 0.56705, 0.56457, 0.56211, 0.55965, 0.5572, 0.55477, 0.55234, 
    0.54993, 0.54752, 0.54512, 0.54274, 0.54036, 0.538, 0.53565, 0.53331, 
    0.53098, 0.52866, 0.52636, 0.52407, 0.52179, 0.51952, 0.51726, 0.51502, 
    0.51279, 0.51057, 0.50836, 0.50616, 0.50397, 0.50179, 0.49962, 0.49746, 
    0.4953, 0.49316, 0.49102, 0.48888, 0.48676, 0.48464, 0.48252, 0.48042, 
    0.47832, 0.47623, 0.47415, 0.47207, 0.47001, 0.46795, 0.46591, 0.46387, 
    0.46185, 0.45984, 0.45783, 0.45584, 0.45386, 0.45188, 0.44992, 0.44797, 
    0.44602, 0.44408, 0.44216, 0.44023, 0.43832, 0.43641, 0.43451, 0.43261, 
    0.43072, 0.42884, 0.42696, 0.42508, 0.42321, 0.42135, 0.41949, 0.41763, 
    0.41579, 0.41394, 0.41211, 0.41027, 0.40845, 0.40663, 0.40482, 0.40301, 
    0.4012, 0.39941, 0.39761, 0.39583, 0.39404, 0.39226, 0.39049, 0.38872, 
    0.38695, 0.38519, 0.38343, 0.38168, 0.37993, 0.37819, 0.37645, 0.37472, 
    0.373, 0.37128, 0.36957, 0.36787, 0.36618, 0.3645, 0.36282, 0.36115, 
    0.35949, 0.35784, 0.3562, 0.35457, 0.35295, 0.35133, 0.34972, 0.34812, 
    0.34652, 0.34493, 0.34335, 0.34177, 0.3402, 0.33863, 0.33707, 0.33552, 
    0.33397, 0.33243, 0.33089, 0.32936, 0.32783, 0.32631, 0.32479, 0.32328, 
    0.32177, 0.32027, 0.31878, 0.31729, 0.31581, 0.31433, 0.31286, 0.3114, 
    0.30994, 0.30848, 0.30703, 0.30559, 0.30416, 0.30272, 0.3013, 0.29988, 
    0.29847, 0.29706, 0.29565, 0.29426, 0.29287, 0.29148, 0.2901, 0.28873, 
    0.28736, 0.286, 0.28465, 0.2833, 0.28196, 0.28062, 0.2793, 0.27797, 
    0.27666, 0.27535, 0.27404, 0.27275, 0.27145, 0.27017, 0.26889, 0.26761, 
    0.26634, 0.26507, 0.26381, 0.26255, 0.26129, 0.26004, 0.25879, 0.25754, 
    0.2563, 0.25506, 0.25381, 0.25257, 0.25134, 0.2501, 0.24887, 0.24764, 
    0.24641, 0.24518, 0.24396, 0.24274, 0.24153, 0.24032, 0.23912, 0.23793, 
    0.23674, 0.23555, 0.23438, 0.23321, 0.23205, 0.2309, 0.22975, 0.22861, 
    0.22748, 0.22636, 0.22525, 0.22414, 0.22304, 0.22194, 0.22085, 0.21977, 
    0.21869, 0.21762, 0.21655, 0.21549, 0.21443, 0.21337, 0.21232, 0.21128, 
    0.21024, 0.2092, 0.20816, 0.20713, 0.20611, 0.20509, 0.20407, 0.20305, 
    0.20204, 0.20104, 0.20003, 0.19904, 0.19804, 0.19705, 0.19607, 0.19509, 
    0.19411, 0.19313, 0.19217, 0.1912, 0.19024, 0.18928, 0.18833, 0.18738, 
    0.18644, 0.18549, 0.18455, 0.18362, 0.18269, 0.18176, 0.18084, 0.17992, 
    0.179, 0.17808, 0.17717, 0.17626, 0.17536, 0.17446, 0.17356, 0.17266, 
    0.17177, 0.17088, 0.16999, 0.16911, 0.16823, 0.16736, 0.16649, 0.16562, 
    0.16476 ;

 press_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 temp =
  267.89, 267.63, 267.36, 267.09, 266.81, 266.53, 266.26, 265.99, 265.72, 
    265.46, 265.2, 264.95, 264.71, 264.49, 264.27, 264.07, 263.88, 263.71, 
    263.55, 263.4, 263.26, 263.14, 263.03, 262.93, 262.84, 262.74, 262.65, 
    262.57, 262.49, 262.42, 262.34, 262.27, 262.21, 262.14, 262.09, 262.04, 
    262, 261.96, 261.93, 261.91, 261.89, 261.87, 261.86, 261.85, 261.85, 
    261.84, 261.84, 261.83, 261.82, 261.82, 261.81, 261.8, 261.79, 261.77, 
    261.76, 261.74, 261.73, 261.71, 261.68, 261.66, 261.64, 261.62, 261.61, 
    261.6, 261.59, 261.58, 261.57, 261.55, 261.54, 261.53, 261.51, 261.5, 
    261.48, 261.46, 261.44, 261.41, 261.39, 261.36, 261.33, 261.3, 261.26, 
    261.23, 261.19, 261.15, 261.12, 261.08, 261.05, 261.02, 260.99, 260.97, 
    260.94, 260.92, 260.89, 260.87, 260.85, 260.84, 260.82, 260.81, 260.79, 
    260.78, 260.77, 260.76, 260.75, 260.74, 260.73, 260.73, 260.72, 260.72, 
    260.71, 260.71, 260.7, 260.7, 260.69, 260.69, 260.69, 260.69, 260.69, 
    260.69, 260.68, 260.68, 260.68, 260.67, 260.66, 260.65, 260.64, 260.63, 
    260.62, 260.6, 260.59, 260.57, 260.55, 260.54, 260.52, 260.51, 260.49, 
    260.47, 260.46, 260.44, 260.43, 260.42, 260.4, 260.39, 260.38, 260.37, 
    260.36, 260.34, 260.33, 260.32, 260.31, 260.29, 260.28, 260.27, 260.26, 
    260.25, 260.23, 260.22, 260.22, 260.21, 260.2, 260.2, 260.19, 260.2, 
    260.2, 260.21, 260.22, 260.23, 260.25, 260.27, 260.29, 260.31, 260.34, 
    260.36, 260.4, 260.43, 260.47, 260.51, 260.55, 260.59, 260.64, 260.69, 
    260.74, 260.8, 260.87, 260.94, 261.02, 261.1, 261.2, 261.31, 261.43, 
    261.56, 261.7, 261.86, 262.02, 262.19, 262.36, 262.53, 262.71, 262.88, 
    263.05, 263.21, 263.38, 263.53, 263.69, 263.85, 264.01, 264.17, 264.34, 
    264.5, 264.67, 264.84, 265.01, 265.17, 265.34, 265.51, 265.68, 265.84, 
    265.99, 266.14, 266.28, 266.42, 266.55, 266.68, 266.8, 266.92, 267.02, 
    267.11, 267.19, 267.26, 267.31, 267.35, 267.38, 267.41, 267.43, 267.45, 
    267.48, 267.5, 267.53, 267.57, 267.61, 267.65, 267.7, 267.75, 267.79, 
    267.83, 267.87, 267.9, 267.93, 267.95, 267.98, 268, 268.01, 268.01, 
    268.01, 268, 268, 268.01, 268.02, 268.02, 268.02, 268.02, 268.02, 268.01, 
    267.99, 267.96, 267.94, 267.92, 267.89, 267.86, 267.82, 267.78, 267.74, 
    267.7, 267.65, 267.59, 267.53, 267.47, 267.41, 267.33, 267.25, 267.17, 
    267.09, 267.01, 266.93, 266.84, 266.75, 266.66, 266.57, 266.48, 266.4, 
    266.31, 266.23, 266.16, 266.08, 266, 265.92, 265.84, 265.77, 265.69, 
    265.62, 265.54, 265.48, 265.43, 265.37, 265.32, 265.28, 265.23, 265.19, 
    265.15, 265.11, 265.07, 265.03, 264.99, 264.96, 264.92, 264.88, 264.84, 
    264.79, 264.75, 264.71, 264.66, 264.62, 264.57, 264.53, 264.49, 264.46, 
    264.42, 264.39, 264.36, 264.33, 264.29, 264.26, 264.22, 264.18, 264.13, 
    264.08, 264.03, 263.98, 263.92, 263.85, 263.78, 263.7, 263.62, 263.54, 
    263.45, 263.37, 263.28, 263.19, 263.11, 263.03, 262.95, 262.87, 262.79, 
    262.72, 262.64, 262.58, 262.51, 262.44, 262.38, 262.32, 262.26, 262.19, 
    262.13, 262.06, 261.99, 261.92, 261.85, 261.78, 261.71, 261.64, 261.58, 
    261.52, 261.46, 261.4, 261.35, 261.3, 261.25, 261.21, 261.17, 261.14, 
    261.11, 261.08, 261.05, 261.02, 260.99, 260.97, 260.94, 260.91, 260.89, 
    260.86, 260.84, 260.81, 260.79, 260.76, 260.74, 260.72, 260.7, 260.68, 
    260.66, 260.65, 260.63, 260.61, 260.59, 260.57, 260.55, 260.53, 260.5, 
    260.48, 260.45, 260.43, 260.4, 260.37, 260.34, 260.31, 260.28, 260.25, 
    260.22, 260.19, 260.16, 260.13, 260.1, 260.07, 260.04, 260.01, 259.98, 
    259.95, 259.92, 259.89, 259.86, 259.82, 259.79, 259.75, 259.72, 259.68, 
    259.65, 259.61, 259.57, 259.54, 259.5, 259.46, 259.43, 259.4, 259.37, 
    259.34, 259.31, 259.28, 259.25, 259.23, 259.2, 259.17, 259.14, 259.11, 
    259.08, 259.05, 259.02, 258.99, 258.95, 258.92, 258.89, 258.86, 258.82, 
    258.79, 258.75, 258.72, 258.69, 258.66, 258.63, 258.6, 258.57, 258.53, 
    258.5, 258.47, 258.44, 258.4, 258.37, 258.33, 258.3, 258.26, 258.22, 
    258.17, 258.13, 258.08, 258.04, 258, 257.96, 257.92, 257.88, 257.84, 
    257.8, 257.77, 257.74, 257.7, 257.68, 257.65, 257.62, 257.59, 257.56, 
    257.54, 257.51, 257.49, 257.46, 257.44, 257.41, 257.38, 257.35, 257.32, 
    257.3, 257.27, 257.24, 257.22, 257.19, 257.17, 257.14, 257.12, 257.09, 
    257.07, 257.05, 257.04, 257.02, 257, 256.98, 256.96, 256.94, 256.93, 
    256.91, 256.89, 256.87, 256.85, 256.83, 256.81, 256.79, 256.77, 256.75, 
    256.73, 256.71, 256.69, 256.67, 256.65, 256.63, 256.61, 256.6, 256.58, 
    256.56, 256.54, 256.52, 256.51, 256.49, 256.47, 256.45, 256.43, 256.41, 
    256.39, 256.37, 256.35, 256.33, 256.31, 256.29, 256.27, 256.25, 256.23, 
    256.21, 256.18, 256.16, 256.14, 256.12, 256.09, 256.07, 256.04, 256.02, 
    256, 255.97, 255.95, 255.93, 255.91, 255.89, 255.87, 255.85, 255.83, 
    255.81, 255.79, 255.78, 255.77, 255.75, 255.74, 255.73, 255.72, 255.71, 
    255.7, 255.69, 255.68, 255.67, 255.66, 255.65, 255.64, 255.63, 255.62, 
    255.61, 255.6, 255.59, 255.58, 255.58, 255.57, 255.56, 255.55, 255.54, 
    255.54, 255.53, 255.52, 255.52, 255.51, 255.5, 255.49, 255.48, 255.46, 
    255.45, 255.43, 255.42, 255.4, 255.38, 255.35, 255.33, 255.31, 255.29, 
    255.27, 255.24, 255.22, 255.19, 255.17, 255.14, 255.12, 255.1, 255.08, 
    255.05, 255.03, 255.01, 254.99, 254.97, 254.95, 254.93, 254.91, 254.89, 
    254.87, 254.85, 254.83, 254.81, 254.79, 254.76, 254.74, 254.71, 254.68, 
    254.66, 254.63, 254.6, 254.58, 254.55, 254.52, 254.49, 254.47, 254.44, 
    254.41, 254.38, 254.35, 254.32, 254.29, 254.27, 254.24, 254.21, 254.18, 
    254.15, 254.13, 254.1, 254.07, 254.04, 254.01, 253.98, 253.95, 253.91, 
    253.88, 253.84, 253.81, 253.77, 253.73, 253.7, 253.66, 253.63, 253.6, 
    253.57, 253.54, 253.51, 253.48, 253.45, 253.43, 253.41, 253.39, 253.38, 
    253.36, 253.35, 253.34, 253.33, 253.32, 253.31, 253.3, 253.29, 253.29, 
    253.28, 253.28, 253.27, 253.27, 253.26, 253.25, 253.24, 253.23, 253.22, 
    253.21, 253.21, 253.2, 253.19, 253.18, 253.17, 253.16, 253.15, 253.15, 
    253.14, 253.13, 253.12, 253.11, 253.1, 253.09, 253.07, 253.06, 253.05, 
    253.03, 253.01, 253, 252.98, 252.96, 252.94, 252.92, 252.9, 252.88, 
    252.86, 252.84, 252.81, 252.79, 252.76, 252.73, 252.71, 252.68, 252.66, 
    252.63, 252.61, 252.58, 252.55, 252.53, 252.5, 252.48, 252.45, 252.43, 
    252.4, 252.37, 252.35, 252.32, 252.29, 252.26, 252.23, 252.2, 252.17, 
    252.14, 252.11, 252.09, 252.06, 252.04, 252.02, 252.01, 252, 251.99, 
    251.99, 251.99, 251.99, 252, 252.01, 252.02, 252.03, 252.05, 252.07, 
    252.09, 252.11, 252.14, 252.17, 252.2, 252.24, 252.28, 252.32, 252.36, 
    252.41, 252.46, 252.52, 252.57, 252.63, 252.7, 252.76, 252.84, 252.91, 
    252.99, 253.07, 253.15, 253.24, 253.33, 253.42, 253.52, 253.62, 253.71, 
    253.81, 253.9, 254, 254.1, 254.2, 254.3, 254.4, 254.5, 254.6, 254.7, 
    254.8, 254.9, 255.01, 255.11, 255.21, 255.31, 255.41, 255.51, 255.6, 
    255.7, 255.79, 255.88, 255.97, 256.06, 256.15, 256.23, 256.31, 256.38, 
    256.46, 256.53, 256.59, 256.65, 256.71, 256.77, 256.81, 256.86, 256.9, 
    256.93, 256.96, 256.99, 257.01, 257.03, 257.04, 257.05, 257.06, 257.06, 
    257.07, 257.07, 257.07, 257.07, 257.07, 257.06, 257.05, 257.04, 257.03, 
    257.01, 257, 256.99, 256.97, 256.95, 256.94, 256.92, 256.91, 256.89, 
    256.88, 256.87, 256.85, 256.84, 256.83, 256.82, 256.81, 256.8, 256.79, 
    256.78, 256.77, 256.76, 256.76, 256.75, 256.74, 256.73, 256.73, 256.72, 
    256.71, 256.7, 256.69, 256.68, 256.67, 256.66, 256.65, 256.64, 256.63, 
    256.62, 256.61, 256.59, 256.58, 256.57, 256.56, 256.55, 256.53, 256.52, 
    256.51, 256.5, 256.48, 256.47, 256.46, 256.44, 256.43, 256.41, 256.4, 
    256.38, 256.36, 256.34, 256.32, 256.3, 256.28, 256.25, 256.23, 256.2, 
    256.18, 256.15, 256.12, 256.09, 256.07, 256.04, 256.01, 255.98, 255.95, 
    255.92, 255.89, 255.86, 255.83, 255.8, 255.77, 255.74, 255.71, 255.68, 
    255.65, 255.62, 255.59, 255.56, 255.53, 255.5, 255.46, 255.43, 255.4, 
    255.36, 255.33, 255.3, 255.26, 255.23, 255.2, 255.17, 255.14, 255.11, 
    255.08, 255.05, 255.02, 254.99, 254.96, 254.93, 254.89, 254.86, 254.83, 
    254.8, 254.76, 254.73, 254.69, 254.66, 254.62, 254.59, 254.55, 254.52, 
    254.48, 254.45, 254.42, 254.38, 254.35, 254.32, 254.29, 254.26, 254.23, 
    254.19, 254.16, 254.13, 254.1, 254.07, 254.04, 254.01, 253.98, 253.95, 
    253.92, 253.89, 253.87, 253.84, 253.81, 253.78, 253.76, 253.73, 253.71, 
    253.68, 253.66, 253.64, 253.62, 253.6, 253.58, 253.56, 253.54, 253.53, 
    253.51, 253.49, 253.48, 253.46, 253.45, 253.44, 253.42, 253.41, 253.39, 
    253.37, 253.36, 253.34, 253.33, 253.31, 253.29, 253.27, 253.26, 253.24, 
    253.22, 253.2, 253.18, 253.16, 253.14, 253.12, 253.1, 253.08, 253.07, 
    253.05, 253.03, 253.01, 252.99, 252.97, 252.95, 252.93, 252.91, 252.89, 
    252.87, 252.84, 252.82, 252.8, 252.77, 252.74, 252.71, 252.68, 252.66, 
    252.63, 252.6, 252.57, 252.54, 252.51, 252.48, 252.45, 252.43, 252.4, 
    252.37, 252.35, 252.32, 252.29, 252.27, 252.24, 252.21, 252.19, 252.16, 
    252.13, 252.1, 252.07, 252.04, 252.01, 251.99, 251.96, 251.93, 251.9, 
    251.87, 251.84, 251.82, 251.79, 251.76, 251.74, 251.71, 251.68, 251.66, 
    251.64, 251.61, 251.59, 251.56, 251.54, 251.52, 251.5, 251.47, 251.45, 
    251.43, 251.41, 251.39, 251.37, 251.35, 251.34, 251.32, 251.3, 251.29, 
    251.27, 251.25, 251.23, 251.22, 251.2, 251.19, 251.17, 251.15, 251.14, 
    251.12, 251.11, 251.09, 251.07, 251.06, 251.04, 251.02, 251, 250.99, 
    250.97, 250.95, 250.93, 250.92, 250.9, 250.88, 250.86, 250.84, 250.82, 
    250.8, 250.77, 250.75, 250.73, 250.7, 250.68, 250.65, 250.62, 250.59, 
    250.56, 250.53, 250.5, 250.47, 250.45, 250.42, 250.39, 250.36, 250.33, 
    250.3, 250.27, 250.24, 250.21, 250.17, 250.14, 250.11, 250.08, 250.05, 
    250.02, 249.98, 249.95, 249.92, 249.88, 249.85, 249.82, 249.79, 249.76, 
    249.72, 249.69, 249.66, 249.63, 249.6, 249.57, 249.54, 249.5, 249.48, 
    249.45, 249.42, 249.39, 249.37, 249.34, 249.32, 249.3, 249.27, 249.25, 
    249.22, 249.2, 249.17, 249.15, 249.12, 249.1, 249.08, 249.05, 249.03, 
    249, 248.98, 248.95, 248.93, 248.91, 248.88, 248.86, 248.84, 248.81, 
    248.79, 248.77, 248.74, 248.72, 248.7, 248.68, 248.66, 248.64, 248.62, 
    248.6, 248.58, 248.56, 248.54, 248.52, 248.5, 248.48, 248.45, 248.43, 
    248.41, 248.39, 248.36, 248.34, 248.31, 248.29, 248.26, 248.24, 248.21, 
    248.19, 248.16, 248.14, 248.11, 248.09, 248.06, 248.04, 248.01, 247.98, 
    247.96, 247.93, 247.91, 247.88, 247.85, 247.83, 247.8, 247.77, 247.74, 
    247.71, 247.68, 247.65, 247.61, 247.58, 247.55, 247.51, 247.48, 247.44, 
    247.41, 247.38, 247.34, 247.31, 247.28, 247.25, 247.22, 247.19, 247.16, 
    247.13, 247.1, 247.08, 247.05, 247.02, 246.99, 246.97, 246.94, 246.91, 
    246.89, 246.87, 246.84, 246.82, 246.8, 246.78, 246.76, 246.74, 246.71, 
    246.69, 246.67, 246.65, 246.63, 246.62, 246.6, 246.58, 246.56, 246.54, 
    246.52, 246.5, 246.48, 246.46, 246.44, 246.42, 246.41, 246.39, 246.37, 
    246.35, 246.33, 246.31, 246.3, 246.28, 246.26, 246.24, 246.23, 246.21, 
    246.19, 246.17, 246.15, 246.13, 246.11, 246.09, 246.07, 246.04, 246.02, 
    246, 245.98, 245.96, 245.94, 245.92, 245.9, 245.88, 245.87, 245.85, 
    245.83, 245.81, 245.79, 245.77, 245.75, 245.73, 245.71, 245.69, 245.67, 
    245.64, 245.62, 245.6, 245.58, 245.56, 245.54, 245.51, 245.49, 245.47, 
    245.45, 245.43, 245.4, 245.38, 245.36, 245.34, 245.32, 245.3, 245.28, 
    245.26, 245.24, 245.22, 245.2, 245.18, 245.16, 245.14, 245.12, 245.1, 
    245.08, 245.06, 245.04, 245.02, 245, 244.98, 244.96, 244.94, 244.92, 
    244.9, 244.89, 244.87, 244.85, 244.84, 244.82, 244.8, 244.79, 244.77, 
    244.75, 244.73, 244.72, 244.7, 244.68, 244.67, 244.65, 244.64, 244.63, 
    244.61, 244.6, 244.58, 244.56, 244.55, 244.53, 244.51, 244.49, 244.47, 
    244.45, 244.43, 244.41, 244.39, 244.37, 244.35, 244.33, 244.31, 244.29, 
    244.27, 244.25, 244.22, 244.2, 244.18, 244.15, 244.13, 244.1, 244.08, 
    244.05, 244.02, 243.99, 243.96, 243.94, 243.91, 243.88, 243.85, 243.82, 
    243.79, 243.75, 243.72, 243.69, 243.66, 243.63, 243.6, 243.57, 243.54, 
    243.51, 243.48, 243.45, 243.42, 243.39, 243.36, 243.33, 243.3, 243.27, 
    243.24, 243.21, 243.18, 243.15, 243.12, 243.09, 243.07, 243.04, 243.01, 
    242.98, 242.96, 242.93, 242.9, 242.87, 242.85, 242.82, 242.8, 242.77, 
    242.75, 242.72, 242.7, 242.67, 242.64, 242.62, 242.59, 242.57, 242.54, 
    242.51, 242.49, 242.46, 242.43, 242.41, 242.38, 242.35, 242.33, 242.3, 
    242.27, 242.25, 242.22, 242.19, 242.17, 242.14, 242.11, 242.09, 242.06, 
    242.03, 242, 241.97, 241.95, 241.92, 241.89, 241.86, 241.83, 241.81, 
    241.78, 241.75, 241.72, 241.7, 241.67, 241.64, 241.62, 241.59, 241.57, 
    241.54, 241.52, 241.49, 241.47, 241.44, 241.42, 241.4, 241.37, 241.35, 
    241.33, 241.3, 241.28, 241.26, 241.24, 241.21, 241.19, 241.17, 241.14, 
    241.12, 241.1, 241.07, 241.05, 241.03, 241.01, 240.98, 240.96, 240.94, 
    240.91, 240.89, 240.86, 240.83, 240.81, 240.78, 240.75, 240.73, 240.7, 
    240.67, 240.64, 240.62, 240.59, 240.56, 240.53, 240.51, 240.48, 240.45, 
    240.42, 240.4, 240.37, 240.34, 240.32, 240.29, 240.26, 240.23, 240.2, 
    240.17, 240.14, 240.11, 240.08, 240.05, 240.02, 239.99, 239.96, 239.93, 
    239.9, 239.87, 239.85, 239.82, 239.79, 239.76, 239.74, 239.71, 239.68, 
    239.65, 239.63, 239.6, 239.57, 239.54, 239.52, 239.49, 239.46, 239.43, 
    239.4, 239.37, 239.34, 239.31, 239.28, 239.25, 239.22, 239.19, 239.16, 
    239.14, 239.11, 239.08, 239.05, 239.02, 238.99, 238.96, 238.94, 238.91, 
    238.88, 238.86, 238.83, 238.8, 238.77, 238.75, 238.72, 238.69, 238.66, 
    238.64, 238.61, 238.58, 238.56, 238.53, 238.5, 238.47, 238.44, 238.41, 
    238.38, 238.36, 238.33, 238.3, 238.27, 238.25, 238.22, 238.19, 238.16, 
    238.13, 238.11, 238.08, 238.05, 238.03, 238, 237.98, 237.95, 237.92, 
    237.9, 237.88, 237.85, 237.83, 237.81, 237.78, 237.76, 237.74, 237.72, 
    237.7, 237.67, 237.65, 237.63, 237.61, 237.59, 237.57, 237.55, 237.53, 
    237.51, 237.49, 237.47, 237.45, 237.43, 237.41, 237.39, 237.37, 237.35, 
    237.33, 237.31, 237.29, 237.27, 237.26, 237.24, 237.22, 237.2, 237.18, 
    237.16, 237.15, 237.13, 237.11, 237.09, 237.07, 237.05, 237.03, 237.01, 
    236.99, 236.96, 236.94, 236.92, 236.9, 236.87, 236.85, 236.82, 236.8, 
    236.77, 236.75, 236.73, 236.7, 236.68, 236.66, 236.63, 236.61, 236.59, 
    236.56, 236.54, 236.51, 236.49, 236.46, 236.44, 236.41, 236.39, 236.36, 
    236.33, 236.3, 236.27, 236.24, 236.21, 236.18, 236.15, 236.13, 236.1, 
    236.07, 236.04, 236.01, 235.98, 235.95, 235.93, 235.9, 235.87, 235.85, 
    235.82, 235.79, 235.77, 235.74, 235.72, 235.69, 235.67, 235.64, 235.61, 
    235.58, 235.55, 235.52, 235.5, 235.47, 235.44, 235.42, 235.39, 235.36, 
    235.34, 235.31, 235.28, 235.26, 235.24, 235.21, 235.19, 235.17, 235.14, 
    235.12, 235.1, 235.07, 235.05, 235.03, 235.01, 234.98, 234.96, 234.93, 
    234.91, 234.88, 234.86, 234.84, 234.81, 234.79, 234.77, 234.74, 234.72, 
    234.7, 234.68, 234.66, 234.64, 234.62, 234.6, 234.58, 234.56, 234.54, 
    234.52, 234.5, 234.48, 234.47, 234.45, 234.43, 234.41, 234.39, 234.38, 
    234.36, 234.34, 234.32, 234.31, 234.29, 234.27, 234.26, 234.24, 234.22, 
    234.21, 234.19, 234.18, 234.16, 234.14, 234.12, 234.1, 234.09, 234.07, 
    234.05, 234.04, 234.02, 234, 233.99, 233.97, 233.95, 233.94, 233.92, 
    233.9, 233.88, 233.86, 233.84, 233.82, 233.8, 233.78, 233.75, 233.73, 
    233.71, 233.68, 233.66, 233.63, 233.6, 233.58, 233.55, 233.53, 233.5, 
    233.47, 233.44, 233.41, 233.38, 233.35, 233.33, 233.3, 233.27, 233.24, 
    233.21, 233.17, 233.14, 233.11, 233.07, 233.04, 233, 232.97, 232.93, 
    232.89, 232.85, 232.81, 232.77, 232.74, 232.7, 232.66, 232.62, 232.59, 
    232.55, 232.51, 232.47, 232.44, 232.4, 232.36, 232.33, 232.29, 232.25, 
    232.22, 232.18, 232.15, 232.11, 232.07, 232.04, 232, 231.97, 231.93, 
    231.9, 231.86, 231.83, 231.79, 231.76, 231.72, 231.69, 231.66, 231.63, 
    231.6, 231.57, 231.54, 231.51, 231.48, 231.45, 231.42, 231.39, 231.36, 
    231.34, 231.31, 231.28, 231.25, 231.22, 231.19, 231.17, 231.14, 231.11, 
    231.08, 231.05, 231.03, 231, 230.97, 230.94, 230.92, 230.89, 230.86, 
    230.84, 230.81, 230.79, 230.76, 230.74, 230.72, 230.69, 230.67, 230.65, 
    230.62, 230.6, 230.58, 230.56, 230.53, 230.51, 230.49, 230.46, 230.44, 
    230.41, 230.39, 230.37, 230.35, 230.33, 230.3, 230.28, 230.26, 230.24, 
    230.22, 230.21, 230.19, 230.17, 230.15, 230.13, 230.11, 230.09, 230.07, 
    230.05, 230.03, 230.01, 229.99, 229.97, 229.94, 229.92, 229.9, 229.88, 
    229.86, 229.84, 229.82, 229.8, 229.78, 229.76, 229.74, 229.72, 229.7, 
    229.69, 229.67, 229.65, 229.63, 229.61, 229.59, 229.58, 229.56, 229.54, 
    229.52, 229.49, 229.47, 229.45, 229.43, 229.4, 229.38, 229.36, 229.33, 
    229.31, 229.29, 229.27, 229.25, 229.23, 229.2, 229.18, 229.16, 229.14, 
    229.12, 229.1, 229.08, 229.06, 229.03, 229.01, 228.99, 228.97, 228.94, 
    228.92, 228.9, 228.88, 228.85, 228.83, 228.8, 228.78, 228.75, 228.73, 
    228.71, 228.68, 228.66, 228.64, 228.61, 228.59, 228.57, 228.55, 228.53, 
    228.51, 228.49, 228.47, 228.45, 228.43, 228.41, 228.39, 228.37, 228.35, 
    228.33, 228.31, 228.29, 228.27, 228.25, 228.23, 228.21, 228.19, 228.16, 
    228.14, 228.12, 228.1, 228.08, 228.05, 228.03, 228.01, 227.99, 227.97, 
    227.95, 227.93, 227.91, 227.89, 227.87, 227.85, 227.83, 227.81, 227.79, 
    227.77, 227.74, 227.72, 227.7, 227.67, 227.65, 227.63, 227.6, 227.58, 
    227.55, 227.53, 227.5, 227.48, 227.45, 227.43, 227.4, 227.38, 227.35, 
    227.33, 227.3, 227.28, 227.26, 227.23, 227.21, 227.19, 227.16, 227.14, 
    227.11, 227.09, 227.06, 227.03, 227.01, 226.98, 226.95, 226.93, 226.9, 
    226.88, 226.85, 226.83, 226.81, 226.78, 226.76, 226.73, 226.71, 226.68, 
    226.66, 226.64, 226.61, 226.58, 226.56, 226.53, 226.51, 226.48, 226.45, 
    226.43, 226.4, 226.38, 226.35, 226.32, 226.29, 226.27, 226.24, 226.21, 
    226.19, 226.16, 226.14, 226.11, 226.09, 226.07, 226.05, 226.02, 226, 
    225.98, 225.96, 225.94, 225.92, 225.9, 225.88, 225.85, 225.83, 225.81, 
    225.79, 225.76, 225.74, 225.72, 225.69, 225.67, 225.65, 225.63, 225.61, 
    225.58, 225.56, 225.54, 225.52, 225.49, 225.47, 225.45, 225.43, 225.41, 
    225.39, 225.37, 225.34, 225.32, 225.3, 225.28, 225.26, 225.24, 225.22, 
    225.2, 225.18, 225.15, 225.13, 225.11, 225.08, 225.05, 225.03, 225, 
    224.98, 224.95, 224.93, 224.91, 224.88, 224.86, 224.83, 224.81, 224.78, 
    224.75, 224.73, 224.7, 224.68, 224.66, 224.63, 224.61, 224.58, 224.56, 
    224.53, 224.51, 224.49, 224.46, 224.44, 224.41, 224.39, 224.36, 224.33, 
    224.31, 224.28, 224.25, 224.22, 224.19, 224.16, 224.13, 224.11, 224.08, 
    224.05, 224.02, 224, 223.97, 223.94, 223.92, 223.89, 223.86, 223.84, 
    223.81, 223.79, 223.76, 223.73, 223.7, 223.68, 223.65, 223.62, 223.59, 
    223.56, 223.53, 223.5, 223.46, 223.43, 223.4, 223.37, 223.34, 223.31, 
    223.28, 223.25, 223.22, 223.19, 223.16, 223.13, 223.1, 223.07, 223.04, 
    223.01, 222.98, 222.95, 222.92, 222.89, 222.86, 222.84, 222.81, 222.78, 
    222.75, 222.72, 222.69, 222.66, 222.63, 222.6, 222.58, 222.55, 222.53, 
    222.51, 222.48, 222.46, 222.43, 222.41, 222.39, 222.37, 222.35, 222.33, 
    222.3, 222.28, 222.25, 222.23, 222.2, 222.18, 222.15, 222.13, 222.1, 
    222.07, 222.04, 222.02, 221.99, 221.97, 221.94, 221.92, 221.89, 221.86, 
    221.83, 221.8, 221.78, 221.75, 221.72, 221.69, 221.66, 221.64, 221.61, 
    221.58, 221.55, 221.52, 221.49, 221.45, 221.42, 221.39, 221.36, 221.33, 
    221.29, 221.26, 221.23, 221.19, 221.16, 221.13, 221.09, 221.06, 221.03, 
    220.99, 220.96, 220.93, 220.9, 220.88, 220.85, 220.82, 220.79, 220.76, 
    220.73, 220.7, 220.68, 220.65, 220.62, 220.6, 220.57, 220.54, 220.52, 
    220.49, 220.46, 220.44, 220.41, 220.39, 220.36, 220.33, 220.31, 220.28, 
    220.26, 220.23, 220.21, 220.19, 220.16, 220.14, 220.12, 220.1, 220.07, 
    220.05, 220.03, 220.01, 219.99, 219.97, 219.95, 219.92, 219.9, 219.88, 
    219.86, 219.84, 219.82, 219.8, 219.78, 219.75, 219.73, 219.71, 219.69, 
    219.67, 219.64, 219.62, 219.6, 219.57, 219.55, 219.52, 219.49, 219.47, 
    219.44, 219.42, 219.39, 219.37, 219.34, 219.32, 219.29, 219.27, 219.24, 
    219.22, 219.19, 219.17, 219.14, 219.11, 219.09, 219.06, 219.04, 219.01, 
    218.99, 218.96, 218.94, 218.91, 218.88, 218.85, 218.82, 218.8, 218.77, 
    218.74, 218.71, 218.68, 218.65, 218.63, 218.6, 218.57, 218.55, 218.52, 
    218.5, 218.47, 218.44, 218.42, 218.39, 218.36, 218.34, 218.31, 218.27, 
    218.24, 218.21, 218.19, 218.16, 218.13, 218.1, 218.07, 218.05, 218.02, 
    217.99, 217.96, 217.93, 217.9, 217.87, 217.85, 217.82, 217.79, 217.76, 
    217.74, 217.71, 217.69, 217.66, 217.64, 217.62, 217.6, 217.57, 217.55, 
    217.53, 217.51, 217.49, 217.47, 217.44, 217.42, 217.4, 217.37, 217.35, 
    217.33, 217.31, 217.29, 217.27, 217.25, 217.23, 217.21, 217.19, 217.17, 
    217.15, 217.13, 217.12, 217.1, 217.08, 217.06, 217.05, 217.03, 217.01, 
    217, 216.98, 216.96, 216.94, 216.92, 216.9, 216.88, 216.86, 216.84, 
    216.81, 216.79, 216.77, 216.75, 216.72, 216.7, 216.68, 216.66, 216.64, 
    216.63, 216.61, 216.59, 216.57, 216.55, 216.53, 216.52, 216.5, 216.47, 
    216.45, 216.43, 216.41, 216.38, 216.36, 216.33, 216.3, 216.28, 216.25, 
    216.22, 216.19, 216.16, 216.13, 216.1, 216.07, 216.05, 216.02, 215.99, 
    215.96, 215.93, 215.91, 215.88, 215.85, 215.82, 215.8, 215.77, 215.74, 
    215.71, 215.68, 215.64, 215.61, 215.58, 215.54, 215.51, 215.48, 215.45, 
    215.42, 215.38, 215.35, 215.32, 215.29, 215.26, 215.23, 215.21, 215.18, 
    215.15, 215.12, 215.09, 215.06, 215.03, 215, 214.97, 214.94, 214.9, 
    214.87, 214.84, 214.81, 214.77, 214.74, 214.71, 214.67, 214.64, 214.61, 
    214.58, 214.55, 214.51, 214.48, 214.45, 214.42, 214.39, 214.36, 214.32, 
    214.29, 214.26, 214.23, 214.2, 214.16, 214.13, 214.1, 214.07, 214.04, 
    214.01, 213.98, 213.95, 213.92, 213.89, 213.86, 213.82, 213.79, 213.76, 
    213.74, 213.71, 213.68, 213.65, 213.62, 213.59, 213.57, 213.54, 213.51, 
    213.48, 213.46, 213.43, 213.4, 213.37, 213.34, 213.32, 213.29, 213.26, 
    213.24, 213.21, 213.19, 213.16, 213.13, 213.11, 213.08, 213.06, 213.03, 
    213, 212.98, 212.95, 212.92, 212.89, 212.87, 212.84, 212.81, 212.79, 
    212.77, 212.74, 212.72, 212.7, 212.67, 212.65, 212.63, 212.61, 212.58, 
    212.56, 212.54, 212.51, 212.49, 212.47, 212.45, 212.43, 212.41, 212.39, 
    212.37, 212.35, 212.33, 212.31, 212.28, 212.26, 212.24, 212.22, 212.2, 
    212.17, 212.15, 212.13, 212.1, 212.08, 212.06, 212.03, 212.01, 211.98, 
    211.96, 211.94, 211.91, 211.89, 211.86, 211.84, 211.81, 211.79, 211.76, 
    211.74, 211.71, 211.69, 211.66, 211.64, 211.61, 211.59, 211.56, 211.54, 
    211.51, 211.49, 211.46, 211.44, 211.42, 211.39, 211.37, 211.34, 211.32, 
    211.3, 211.28, 211.25, 211.23, 211.21, 211.19, 211.17, 211.15, 211.12, 
    211.1, 211.08, 211.06, 211.04, 211.02, 211, 210.97, 210.95, 210.93, 
    210.91, 210.89, 210.86, 210.84, 210.82, 210.8, 210.78, 210.75, 210.73, 
    210.71, 210.69, 210.67, 210.65, 210.63, 210.61, 210.59, 210.57, 210.54, 
    210.52, 210.5, 210.48, 210.46, 210.44, 210.42, 210.4, 210.38, 210.36, 
    210.34, 210.32, 210.3, 210.28, 210.26, 210.24, 210.22, 210.21, 210.19, 
    210.17, 210.15, 210.13, 210.12, 210.1, 210.08, 210.06, 210.04, 210.02, 
    209.99, 209.97, 209.95, 209.92, 209.9, 209.87, 209.85, 209.82, 209.8, 
    209.77, 209.75, 209.72, 209.7, 209.68, 209.66, 209.63, 209.61, 209.59, 
    209.57, 209.54, 209.52, 209.5, 209.47, 209.45, 209.43, 209.4, 209.38, 
    209.35, 209.32, 209.3, 209.27, 209.24, 209.22, 209.19, 209.16, 209.13, 
    209.11, 209.08, 209.05, 209.03, 209, 208.98, 208.96, 208.93, 208.91, 
    208.88, 208.86, 208.84, 208.81, 208.78, 208.76, 208.73, 208.7, 208.67, 
    208.64, 208.62, 208.59, 208.56, 208.54, 208.51, 208.48, 208.45, 208.43, 
    208.4, 208.38, 208.35, 208.32, 208.3, 208.27, 208.24, 208.21, 208.18, 
    208.15, 208.13, 208.1, 208.08, 208.05, 208.03, 208, 207.98, 207.95, 
    207.93, 207.91, 207.88, 207.86, 207.84, 207.81, 207.79, 207.76, 207.74, 
    207.71, 207.69, 207.66, 207.64, 207.61, 207.59, 207.56, 207.53, 207.51, 
    207.48, 207.45, 207.43, 207.4, 207.38, 207.35, 207.33, 207.31, 207.29, 
    207.27, 207.25, 207.23, 207.21, 207.19, 207.17, 207.14, 207.12, 207.1, 
    207.07, 207.05, 207.02, 207, 206.97, 206.95, 206.92, 206.9, 206.87, 
    206.85, 206.82, 206.8, 206.77, 206.74, 206.72, 206.69, 206.67, 206.65, 
    206.62, 206.6, 206.57, 206.55, 206.52, 206.5, 206.47, 206.45, 206.42, 
    206.4, 206.37, 206.34, 206.32, 206.29, 206.26, 206.24, 206.21, 206.18, 
    206.15, 206.13, 206.1, 206.08, 206.05, 206.03, 206.01, 205.98, 205.96, 
    205.93, 205.91, 205.89, 205.87, 205.85, 205.83, 205.8, 205.78, 205.76, 
    205.73, 205.71, 205.68, 205.66, 205.64, 205.62, 205.59, 205.57, 205.55, 
    205.52, 205.5, 205.48, 205.45, 205.43, 205.4, 205.38, 205.35, 205.32, 
    205.3, 205.27, 205.24, 205.21, 205.19, 205.16, 205.13, 205.1, 205.07, 
    205.04, 205.01, 204.98, 204.95, 204.92, 204.89, 204.86, 204.83, 204.8, 
    204.77, 204.74, 204.71, 204.68, 204.65, 204.61, 204.58, 204.55, 204.52, 
    204.49, 204.46, 204.42, 204.4, 204.37, 204.34, 204.31, 204.29, 204.27, 
    204.24, 204.22, 204.19, 204.17, 204.15, 204.12, 204.1, 204.07, 204.05, 
    204.03, 204.01, 203.98, 203.96, 203.94, 203.91, 203.89, 203.87, 203.85, 
    203.83, 203.81, 203.79, 203.78, 203.76, 203.74, 203.73, 203.71, 203.7, 
    203.68, 203.67, 203.66, 203.64, 203.63, 203.62, 203.6, 203.59, 203.57, 
    203.56, 203.55, 203.53, 203.52, 203.51, 203.5, 203.49, 203.48, 203.47, 
    203.46, 203.44, 203.43, 203.42, 203.41, 203.41, 203.4, 203.39, 203.39, 
    203.38, 203.37, 203.37, 203.37, 203.36, 203.36, 203.35, 203.35, 203.35, 
    203.34, 203.34, 203.33, 203.32, 203.31, 203.31, 203.3, 203.29, 203.29, 
    203.29, 203.28, 203.28, 203.27, 203.27, 203.27, 203.26, 203.26, 203.26, 
    203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 203.26, 
    203.26, 203.26, 203.25, 203.25, 203.24, 203.24, 203.23, 203.23, 203.23, 
    203.22, 203.22, 203.22, 203.23, 203.23, 203.23, 203.24, 203.24, 203.24, 
    203.25, 203.25, 203.25, 203.26, 203.26, 203.27, 203.27, 203.27, 203.28, 
    203.28, 203.29, 203.3, 203.3, 203.31, 203.32, 203.32, 203.33, 203.34, 
    203.35, 203.36, 203.37, 203.38, 203.39, 203.4, 203.41, 203.43, 203.44, 
    203.45, 203.46, 203.47, 203.48, 203.5, 203.51, 203.52, 203.54, 203.55, 
    203.56, 203.58, 203.59, 203.61, 203.62, 203.64, 203.65, 203.66, 203.68, 
    203.69, 203.7, 203.71, 203.72, 203.73, 203.75, 203.76, 203.78, 203.79, 
    203.81, 203.83, 203.84, 203.86, 203.88, 203.9, 203.93, 203.95, 203.97, 
    204, 204.02, 204.04, 204.06, 204.09, 204.11, 204.13, 204.15, 204.17, 
    204.19, 204.21, 204.23, 204.24, 204.25, 204.26, 204.28, 204.29, 204.3, 
    204.31, 204.32, 204.33, 204.34, 204.34, 204.35, 204.36, 204.36, 204.36, 
    204.36, 204.35, 204.35, 204.34, 204.33, 204.32, 204.31, 204.3, 204.29, 
    204.27, 204.26, 204.24, 204.23, 204.21, 204.19, 204.17, 204.15, 204.13, 
    204.11, 204.08, 204.06, 204.04, 204.02, 204, 203.98, 203.96, 203.94, 
    203.92, 203.9, 203.88, 203.86, 203.84, 203.83, 203.81, 203.79, 203.78, 
    203.76, 203.75, 203.74, 203.73, 203.71, 203.7, 203.69, 203.67, 203.66, 
    203.65, 203.63, 203.61, 203.6, 203.58, 203.56, 203.54, 203.52, 203.5, 
    203.48, 203.47, 203.45, 203.43, 203.41, 203.39, 203.37, 203.35, 203.34, 
    203.32, 203.3, 203.28, 203.26, 203.24, 203.22, 203.2, 203.18, 203.17, 
    203.14, 203.12, 203.1, 203.08, 203.06, 203.03, 203.01, 202.99, 202.97, 
    202.95, 202.93, 202.91, 202.89, 202.88, 202.86, 202.85, 202.83, 202.82, 
    202.81, 202.79, 202.78, 202.78, 202.77, 202.76, 202.76, 202.75, 202.75, 
    202.75, 202.75, 202.75, 202.76, 202.76, 202.77, 202.78, 202.79, 202.8, 
    202.81, 202.81, 202.82, 202.83, 202.84, 202.85, 202.86, 202.87, 202.87, 
    202.88, 202.89, 202.9, 202.91, 202.92, 202.93, 202.94, 202.95, 202.96, 
    202.97, 202.98, 202.99, 203, 203.01, 203.02, 203.03, 203.04, 203.04, 
    203.05, 203.06, 203.06, 203.07, 203.07, 203.08, 203.08, 203.08, 203.09, 
    203.09, 203.09, 203.1, 203.1, 203.11, 203.11, 203.12, 203.12, 203.13, 
    203.14, 203.15, 203.16, 203.17, 203.19, 203.2, 203.22, 203.24, 203.26, 
    203.28, 203.3, 203.32, 203.34, 203.36, 203.38, 203.39, 203.41, 203.43, 
    203.45, 203.46, 203.47, 203.49, 203.5, 203.51, 203.51, 203.52, 203.53, 
    203.55, 203.56, 203.57, 203.58, 203.59, 203.6, 203.61, 203.62, 203.63, 
    203.63, 203.64, 203.65, 203.65, 203.66, 203.66, 203.66, 203.65, 203.65, 
    203.64, 203.64, 203.63, 203.63, 203.63, 203.63, 203.63, 203.63, 203.64, 
    203.64, 203.65, 203.66, 203.67, 203.69, 203.7, 203.72, 203.73, 203.75, 
    203.77, 203.79, 203.8, 203.82, 203.83, 203.85, 203.87, 203.89, 203.91, 
    203.92, 203.94, 203.96, 203.98, 204, 204.03, 204.05, 204.07, 204.09, 
    204.12, 204.14, 204.16, 204.18, 204.2, 204.21, 204.23, 204.25, 204.26, 
    204.27, 204.29, 204.3, 204.31, 204.33, 204.34, 204.36, 204.37, 204.39, 
    204.4, 204.42, 204.43, 204.45, 204.46, 204.48, 204.49, 204.51, 204.53, 
    204.54, 204.56, 204.57, 204.59, 204.61, 204.63, 204.65, 204.67, 204.69, 
    204.71, 204.73, 204.75, 204.78, 204.8, 204.83, 204.86, 204.88, 204.91, 
    204.94, 204.96, 204.99, 205.01, 205.03, 205.05, 205.07, 205.08, 205.09, 
    205.11, 205.12, 205.13, 205.14, 205.15, 205.17, 205.18, 205.19, 205.21, 
    205.22, 205.23, 205.25, 205.26, 205.28, 205.29, 205.31, 205.32, 205.33, 
    205.35, 205.36, 205.38, 205.39, 205.4, 205.42, 205.43, 205.45, 205.46, 
    205.47, 205.49, 205.5, 205.51, 205.52, 205.53, 205.54, 205.55, 205.56, 
    205.57, 205.58, 205.59, 205.6, 205.61, 205.62, 205.63, 205.63, 205.64, 
    205.64, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 205.65, 
    205.65, 205.65, 205.64, 205.64, 205.63, 205.62, 205.61, 205.6, 205.58, 
    205.57, 205.56, 205.55, 205.54, 205.53, 205.51, 205.5, 205.49, 205.49, 
    205.48, 205.48, 205.48, 205.48, 205.47, 205.47, 205.48, 205.48, 205.48, 
    205.49, 205.5, 205.51, 205.52, 205.53, 205.54, 205.55, 205.55, 205.56, 
    205.57, 205.58, 205.59, 205.59, 205.6, 205.61, 205.62, 205.63, 205.64, 
    205.65, 205.66, 205.68, 205.69, 205.7, 205.72, 205.73, 205.75, 205.77, 
    205.78, 205.8, 205.81, 205.82, 205.84, 205.85, 205.87, 205.88, 205.89, 
    205.91, 205.92, 205.93, 205.94, 205.94, 205.95, 205.96, 205.97, 205.98, 
    205.99, 206, 206.01, 206.02, 206.04, 206.05, 206.07, 206.08, 206.1, 
    206.12, 206.13, 206.15, 206.17, 206.19, 206.21, 206.23, 206.25, 206.26, 
    206.28, 206.3, 206.31, 206.33, 206.34, 206.36, 206.37, 206.39, 206.4, 
    206.41, 206.43, 206.44, 206.45, 206.46, 206.47, 206.48, 206.49, 206.49, 
    206.5, 206.5, 206.5, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 
    206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 206.51, 
    206.51, 206.51, 206.52, 206.52, 206.52, 206.52, 206.52, 206.52, 206.53, 
    206.53, 206.53, 206.53, 206.53, 206.53, 206.54, 206.54, 206.54, 206.54, 
    206.55, 206.55, 206.56, 206.57, 206.58, 206.59, 206.6, 206.61, 206.62, 
    206.63, 206.64, 206.66, 206.67, 206.68, 206.69, 206.7, 206.71, 206.71, 
    206.72, 206.73, 206.73, 206.74, 206.75, 206.76, 206.77, 206.78, 206.79, 
    206.8, 206.81, 206.83, 206.84, 206.85, 206.87, 206.88, 206.89, 206.9, 
    206.91, 206.92, 206.93, 206.94, 206.95, 206.96, 206.97, 206.98, 206.99, 
    207, 207, 207.01, 207.02, 207.03, 207.03, 207.04, 207.04, 207.05, 207.05, 
    207.06, 207.06, 207.07, 207.07, 207.07, 207.07, 207.08, 207.08, 207.07, 
    207.07, 207.07, 207.06, 207.06, 207.06, 207.05, 207.05, 207.04, 207.04, 
    207.03, 207.03, 207.03, 207.02, 207.02, 207.02, 207.02, 207.02, 207.02, 
    207.02, 207.01, 207.01, 207, 207, 206.99, 206.98, 206.97, 206.95, 206.96, 
    206.97, 206.98, 206.99, 207, 207.01, 207.02, 207.03, 207.04, 207.04, 
    207.05, 207.05, 207.06, 207.06, 207.06, 207.06, 207.06, 207.05, 207.05, 
    207.04, 207.03, 207.02, 207.01, 207, 206.99, 206.97, 206.96, 206.95, 
    206.94, 206.92, 206.91, 206.9, 206.9, 206.89, 206.88, 206.88, 206.87, 
    206.87, 206.87, 206.86, 206.86, 206.86, 206.86, 206.86, 206.86, 206.86, 
    206.86, 206.86, 206.86, 206.85, 206.85, 206.85, 206.85, 206.84, 206.84, 
    206.84, 206.83, 206.83, 206.82, 206.82, 206.81, 206.81, 206.81, 206.8, 
    206.8, 206.8, 206.79, 206.79, 206.79, 206.79, 206.79, 206.79, 206.8, 
    206.8, 206.8, 206.8, 206.81, 206.81, 206.81, 206.82, 206.82, 206.82, 
    206.82, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 206.83, 
    206.83, 206.83, 206.83, 206.82, 206.82, 206.82, 206.82, 206.81, 206.81, 
    206.81, 206.8, 206.8, 206.8, 206.8, 206.79, 206.79, 206.79, 206.78, 
    206.78, 206.78, 206.78, 206.77, 206.77, 206.77, 206.77, 206.77, 206.76, 
    206.76, 206.76, 206.76, 206.76, 206.75, 206.75, 206.75, 206.75, 206.74, 
    206.74, 206.74, 206.73, 206.73, 206.73, 206.72, 206.72, 206.71, 206.7, 
    206.69, 206.69, 206.68, 206.67, 206.65, 206.64, 206.63, 206.61, 206.6, 
    206.58, 206.56, 206.54, 206.52, 206.49, 206.47, 206.44, 206.41, 206.39, 
    206.36, 206.32, 206.29, 206.26, 206.23, 206.19, 206.16, 206.12, 206.09, 
    206.05, 206.02, 205.98, 205.94, 205.91, 205.87, 205.83, 205.8, 205.76, 
    205.73, 205.69, 205.65, 205.62, 205.58, 205.55, 205.51, 205.48, 205.44, 
    205.41, 205.37, 205.33, 205.3, 205.26, 205.23, 205.19, 205.16, 205.12, 
    205.08, 205.05, 205.01, 204.97, 204.93, 204.89, 204.86, 204.82, 204.77, 
    204.73, 204.69, 204.65, 204.6, 204.55, 204.5, 204.45, 204.4, 204.35, 
    204.29, 204.23, 204.17, 204.11, 204.05, 203.98, 203.91, 203.84, 203.77, 
    203.7, 203.62, 203.55, 203.47, 203.4, 203.32, 203.25, 203.17, 203.1, 
    203.03, 202.96, 202.89, 202.82, 202.75, 202.69, 202.63, 202.57, 202.51, 
    202.45, 202.4, 202.35, 202.3, 202.25, 202.21, 202.16, 202.12, 202.08, 
    202.05, 202.01, 201.98, 201.95, 201.93, 201.9, 201.88, 201.87, 201.85, 
    201.84, 201.83, 201.82, 201.82, 201.82, 201.82, 201.82, 201.83, 201.84, 
    201.85, 201.86, 201.87, 201.88, 201.9, 201.91, 201.93, 201.95, 201.96, 
    201.98, 201.99, 202.01, 202.02, 202.04, 202.05, 202.06, 202.07, 202.08, 
    202.09, 202.09, 202.1, 202.1, 202.1, 202.1, 202.1, 202.1, 202.1, 202.09, 
    202.09, 202.08, 202.07, 202.06, 202.05, 202.04, 202.03, 202.01, 201.99, 
    201.97, 201.95, 201.93, 201.9, 201.87, 201.84, 201.81, 201.77, 201.73, 
    201.69, 201.65, 201.6, 201.55, 201.5, 201.44, 201.39, 201.33, 201.27, 
    201.2, 201.14, 201.07, 201.01, 200.94, 200.87, 200.8, 200.73, 200.65, 
    200.58, 200.51, 200.44, 200.37, 200.29, 200.22, 200.15, 200.09, 200.02, 
    199.95, 199.89, 199.83, 199.77, 199.71, 199.65, 199.6, 199.55, 199.5, 
    199.46, 199.42, 199.38, 199.34, 199.31, 199.28, 199.25, 199.23, 199.21, 
    199.19, 199.18, 199.16, 199.15, 199.15, 199.14, 199.14, 199.14, 199.15, 
    199.15, 199.16, 199.17, 199.18, 199.19, 199.21, 199.22, 199.24, 199.26, 
    199.28, 199.3, 199.32, 199.35, 199.37, 199.39, 199.42, 199.44, 199.47, 
    199.49, 199.52, 199.55, 199.57, 199.6, 199.62, 199.65, 199.67, 199.7, 
    199.72, 199.75, 199.77, 199.8, 199.82, 199.84, 199.86, 199.88, 199.9, 
    199.91, 199.93, 199.94, 199.95, 199.96, 199.97, 199.98, 199.98, 199.98, 
    199.98, 199.98, 199.98, 199.97, 199.97, 199.96, 199.96, 199.95, 199.94, 
    199.93, 199.93, 199.92, 199.91, 199.91, 199.91, 199.9, 199.9, 199.9, 
    199.9, 199.9, 199.91, 199.91, 199.92, 199.92, 199.93, 199.94, 199.95, 
    199.96, 199.97, 199.98, 199.98, 199.99, 200, 200.01, 200.01, 200.02, 
    200.03, 200.03, 200.03, 200.04, 200.04, 200.04, 200.04, 200.04, 200.04, 
    200.04, 200.04, 200.04, 200.03, 200.03, 200.02, 200.01, 200, 199.99, 
    199.98, 199.96, 199.95, 199.93, 199.91, 199.88, 199.86, 199.83, 199.81, 
    199.78, 199.75, 199.72, 199.69, 199.66, 199.63, 199.6, 199.57, 199.54, 
    199.52, 199.49, 199.47, 199.46, 199.44, 199.43, 199.43, 199.42, 199.42, 
    199.43, 199.44, 199.45, 199.47, 199.49, 199.52, 199.54, 199.58, 199.61, 
    199.65, 199.69, 199.73, 199.78, 199.82, 199.87, 199.92, 199.96, 200.01, 
    200.06, 200.1, 200.14, 200.18, 200.22, 200.26, 200.29, 200.31, 200.33, 
    200.35, 200.36, 200.37, 200.37, 200.37, 200.36, 200.35, 200.33, 200.31, 
    200.28, 200.25, 200.21, 200.17, 200.13, 200.09, 200.04, 199.99, 199.94, 
    199.89, 199.84, 199.8, 199.75, 199.7, 199.66, 199.62, 199.58, 199.54, 
    199.51, 199.48, 199.45, 199.43, 199.4, 199.39, 199.37, 199.36, 199.35, 
    199.34, 199.34, 199.34, 199.34, 199.35, 199.35, 199.36, 199.38, 199.4, 
    199.42, 199.44, 199.47, 199.5, 199.54, 199.58, 199.62, 199.67, 199.72, 
    199.78, 199.84, 199.91, 199.97, 200.04, 200.12, 200.19, 200.26, 200.34, 
    200.42, 200.49, 200.57, 200.64, 200.72, 200.79, 200.85, 200.92, 200.98, 
    201.04, 201.09, 201.14, 201.18, 201.22, 201.26, 201.29, 201.31, 201.33, 
    201.35, 201.36, 201.37, 201.37, 201.36, 201.36, 201.34, 201.33, 201.3, 
    201.28, 201.25, 201.22, 201.19, 201.15, 201.11, 201.07, 201.03, 200.99, 
    200.95, 200.91, 200.88, 200.84, 200.81, 200.78, 200.75, 200.73, 200.7, 
    200.69, 200.67, 200.66, 200.66, 200.65, 200.66, 200.66, 200.67, 200.68, 
    200.69, 200.71, 200.73, 200.76, 200.79, 200.82, 200.86, 200.9, 200.94, 
    200.99, 201.04, 201.09, 201.15, 201.21, 201.27, 201.33, 201.39, 201.46, 
    201.53, 201.6, 201.67, 201.75, 201.83, 201.9, 201.98, 202.07, 202.15, 
    202.24, 202.33, 202.42, 202.52, 202.61, 202.71, 202.82, 202.92, 203.02, 
    203.13, 203.23, 203.34, 203.44, 203.54, 203.64, 203.73, 203.82, 203.9, 
    203.98, 204.05, 204.11, 204.17, 204.22, 204.26, 204.29, 204.31, 204.33, 
    204.33, 204.33, 204.32, 204.3, 204.27, 204.24, 204.2, 204.15, 204.09, 
    204.03, 203.97, 203.9, 203.83, 203.75, 203.68, 203.6, 203.53, 203.45, 
    203.38, 203.32, 203.26, 203.2, 203.15, 203.11, 203.08, 203.06, 203.04, 
    203.03, 203.04, 203.05, 203.07, 203.1, 203.14, 203.18, 203.24, 203.3, 
    203.37, 203.45, 203.53, 203.62, 203.71, 203.81, 203.92, 204.03, 204.14, 
    204.26, 204.38, 204.5, 204.63, 204.76, 204.89, 205.02, 205.16, 205.29, 
    205.43, 205.57, 205.71, 205.86, 206, 206.15, 206.29, 206.44, 206.59, 
    206.74, 206.9, 207.05, 207.21, 207.36, 207.52, 207.68, 207.85, 208.01, 
    208.18, 208.35, 208.52, 208.69, 208.87, 209.05, 209.23, 209.41, 209.59, 
    209.77, 209.96, 210.15, 210.33, 210.52, 210.71, 210.9, 211.08, 211.26, 
    211.44, 211.62, 211.8, 211.96, 212.13, 212.29, 212.44, 212.58, 212.72, 
    212.84, 212.96, 213.08, 213.18, 213.28, 213.36, 213.44, 213.51, 213.58, 
    213.64, 213.69, 213.74, 213.79, 213.84, 213.88, 213.92, 213.96, 214.01, 
    214.05, 214.1, 214.15, 214.21, 214.27, 214.33, 214.4, 214.47, 214.55, 
    214.63, 214.72, 214.81, 214.91, 215.01, 215.11, 215.22, 215.33, 215.45, 
    215.56, 215.68, 215.79, 215.91, 216.03, 216.14, 216.26, 216.37, 216.48, 
    216.59, 216.69, 216.79, 216.88, 216.98, 217.06, 217.14, 217.22, 217.3, 
    217.36, 217.43, 217.49, 217.55, 217.61, 217.66, 217.72, 217.77, 217.82, 
    217.88, 217.93, 217.98, 218.04, 218.1, 218.16, 218.22, 218.28, 218.34, 
    218.41, 218.47, 218.54, 218.61, 218.68, 218.74, 218.81, 218.88, 218.94, 
    219.01, 219.07, 219.14, 219.2, 219.26, 219.33, 219.39, 219.45, 219.52, 
    219.58, 219.65, 219.72, 219.79, 219.87, 219.95, 220.04, 220.13, 220.23, 
    220.33, 220.44, 220.55, 220.67, 220.8, 220.94, 221.09, 221.24, 221.4, 
    221.56, 221.74, 221.92, 222.1, 222.29, 222.49, 222.69, 222.89, 223.1, 
    223.31, 223.53, 223.74, 223.96, 224.18, 224.4, 224.62, 224.84, 225.06, 
    225.28, 225.5, 225.71, 225.93, 226.14, 226.35, 226.56, 226.77, 226.97, 
    227.17, 227.36, 227.55, 227.74, 227.92, 228.1, 228.27, 228.43, 228.6, 
    228.75, 228.91, 229.06, 229.2, 229.35, 229.49, 229.63, 229.77, 229.91, 
    230.05, 230.2, 230.35, 230.5, 230.65, 230.81, 230.97, 231.13, 231.3, 
    231.47, 231.64, 231.81, 231.98, 232.15, 232.32, 232.48, 232.64, 232.8, 
    232.95, 233.09, 233.23, 233.37, 233.5, 233.62, 233.74, 233.85, 233.97, 
    234.07, 234.18, 234.28, 234.39, 234.49, 234.6, 234.71, 234.82, 234.94, 
    235.06, 235.19, 235.33, 235.47, 235.62, 235.78, 235.95, 236.13, 236.32, 
    236.51, 236.72, 236.93, 237.15, 237.38, 237.61, 237.86, 238.11, 238.36, 
    238.62, 238.88, 239.15, 239.42, 239.69, 239.96, 240.24, 240.5, 240.77, 
    241.04, 241.3, 241.55, 241.8, 242.05, 242.28, 242.51, 242.73, 242.95, 
    243.15, 243.34, 243.53, 243.71, 243.87, 244.03, 244.18, 244.33, 244.46, 
    244.59, 244.71, 244.82, 244.93, 245.03, 245.13, 245.23, 245.32, 245.42, 
    245.51, 245.61, 245.71, 245.81, 245.91, 246.02, 246.13, 246.25, 246.37, 
    246.5, 246.64, 246.78, 246.93, 247.09, 247.25, 247.42, 247.6, 247.78, 
    247.96, 248.15, 248.35, 248.55, 248.75, 248.96, 249.17, 249.38, 249.6, 
    249.82, 250.04, 250.26, 250.49, 250.72, 250.95, 251.18, 251.42, 251.65, 
    251.89, 252.13, 252.36, 252.6, 252.84, 253.07, 253.31, 253.55, 253.78, 
    254.01, 254.25, 254.48, 254.71, 254.93, 255.16, 255.38, 255.61, 255.83, 
    256.05, 256.27, 256.49, 256.71, 256.92, 257.14, 257.36, 257.57, 257.79, 
    258, 258.21, 258.43, 258.64, 258.85, 259.06, 259.27, 259.48, 259.69, 
    259.9, 260.11, 260.32, 260.52, 260.73, 260.94, 261.14, 261.35, 261.56, 
    261.77, 261.98, 262.19, 262.4, 262.61, 262.83, 263.04, 263.26, 263.48, 
    263.7, 263.92, 264.14, 264.36, 264.59, 264.81, 265.04, 265.26, 265.49, 
    265.72, 265.95, 266.17, 266.4, 266.63, 266.86, 267.09, 267.32, 267.55, 
    267.77, 268, 268.22, 268.45, 268.67, 268.89, 269.11, 269.32, 269.53, 
    269.75, 269.95, 270.16, 270.36, 270.56, 270.76, 270.96, 271.15, 271.34, 
    271.53, 271.71, 271.9, 272.08, 272.26, 272.44, 272.62, 272.8, 272.98, 
    273.16, 273.33, 273.51, 273.68, 273.86, 274.04, 274.21, 274.39, 274.57, 
    274.74, 274.92, 275.1, 275.27, 275.45, 275.63, 275.81, 275.99, 276.17, 
    276.35, 276.52, 276.7, 276.88, 277.06, 277.23, 277.41, 277.58, 277.75, 
    277.92, 278.08, 278.25, 278.41, 278.57, 278.72, 278.88, 279.03, 279.18, 
    279.32, 279.47, 279.61, 279.75, 279.9, 280.04, 280.18, 280.33, 280.48, 
    280.63, 280.79, 280.95, 281.11, 281.28, 281.45, 281.63, 281.81, 281.99, 
    282.18, 282.37, 282.57, 282.76, 282.96, 283.16, 283.36, 283.55, 283.75, 
    283.94, 284.13, 284.32, 284.5, 284.68, 284.86, 285.02, 285.19, 285.35, 
    285.5, 285.65, 285.79, 285.92, 286.05, 286.18, 286.3, 286.41, 286.52, 
    286.62, 286.72, 286.82, 286.91, 287, 287.09, 287.18, 287.26, 287.35, 
    287.43, 287.51, 287.6, 287.68, 287.77, 287.86, 287.95, 288.04, 288.14, 
    288.24, 288.33, 288.44, 288.54, 288.65, 288.75, 288.86, 288.97, 289.09, 
    289.2, 289.31, 289.42, 289.53, 289.65, 289.76, 289.86, 289.97, 290.07, 
    290.17, 290.27, 290.37, 290.46, 290.55, 290.63, 290.71, 290.78, 290.85, 
    290.92, 290.98, 291.04, 291.09, 291.14, 291.18, 291.22, 291.25, 291.28, 
    291.31, 291.33, 291.34, 291.35, 291.35, 291.35, 291.34, 291.32, 291.3, 
    291.27, 291.23, 291.19, 291.14, 291.08, 291.01, 290.93, 290.83, 290.72, 
    290.59, 290.46, 290.33, 290.19, 290.05, 289.91, 289.77, 289.62, 289.48, 
    289.34, 289.19, 289.05, 288.91, 288.76, 288.62, 288.48, 288.34, 288.2, 
    288.06, 287.92, 287.79, 287.65, 287.51, 287.38, 287.24, 287.11, 286.97, 
    286.84, 286.7, 286.57, 286.43, 286.3, 286.16, 286.02, 285.89, 285.75, 
    285.62, 285.48, 285.34, 285.21, 285.07, 284.93, 284.8, 284.66, 284.53, 
    284.39, 284.26, 284.12, 283.99, 283.85, 283.72, 283.58, 283.45, 283.31, 
    283.17, 283.03, 282.9, 282.76, 282.62, 282.47, 282.33, 282.19, 282.04, 
    281.9, 281.75, 281.6, 281.45, 281.3, 281.15, 281, 280.85, 280.7, 280.55, 
    280.39, 280.24, 280.09, 279.94, 279.79, 279.63, 279.48, 279.33, 279.17, 
    279.02, 278.86, 278.71, 278.55, 278.39, 278.23, 278.07, 277.91, 277.74, 
    277.58, 277.41, 277.24, 277.08, 276.91, 276.73, 276.56, 276.39, 276.22, 
    276.04, 275.87, 275.69, 275.51, 275.33, 275.15, 274.97, 274.79, 274.61, 
    274.43, 274.24, 274.06, 273.87, 273.69, 273.5, 273.31, 273.12, 272.93, 
    272.74, 272.55, 272.35, 272.16, 271.97, 271.78, 271.59, 271.4, 271.2, 
    271.01, 270.82, 270.64, 270.45, 270.26, 270.07, 269.88, 269.7, 269.51, 
    269.32, 269.13, 268.95, 268.76, 268.57, 268.38, 268.19, 268, 267.81, 
    267.62, 267.43, 267.24, 267.05, 266.85, 266.66, 266.47, 266.27, 266.08, 
    265.88, 265.69, 265.49, 265.29, 265.1, 264.9, 264.7, 264.5, 264.31, 
    264.11, 263.91, 263.71, 263.51, 263.31, 263.11, 262.91, 262.71, 262.51, 
    262.3, 262.1, 261.9, 261.7, 261.5, 261.29, 261.09, 260.89, 260.69, 
    260.48, 260.28, 260.08, 259.87, 259.67, 259.47, 259.26, 259.06, 258.86, 
    258.65, 258.45, 258.25, 258.04, 257.84, 257.63, 257.42, 257.22, 257.01, 
    256.8, 256.59, 256.38, 256.16, 255.95, 255.74, 255.52, 255.3, 255.09, 
    254.87, 254.65, 254.43, 254.21, 253.99, 253.77, 253.55, 253.34, 253.12, 
    252.9, 252.69, 252.47, 252.26, 252.05, 251.84, 251.63, 251.43, 251.22, 
    251.02, 250.82, 250.61, 250.41, 250.22, 250.02, 249.82, 249.62, 249.43, 
    249.23, 249.04, 248.84, 248.65, 248.46, 248.26, 248.07, 247.88, 247.68, 
    247.49, 247.3, 247.11, 246.92, 246.73, 246.54, 246.35, 246.16, 245.97, 
    245.78, 245.59, 245.41, 245.22, 245.04, 244.85, 244.67, 244.49, 244.31, 
    244.13, 243.95, 243.77, 243.59, 243.41, 243.24, 243.06, 242.89, 242.72, 
    242.55, 242.38, 242.21, 242.05, 241.88, 241.72, 241.56, 241.4, 241.24, 
    241.09, 240.94, 240.79, 240.64, 240.5, 240.36, 240.23, 240.1, 239.97, 
    239.85, 239.74, 239.63 ;

 temp_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 shum =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 shum_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 meteo_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;
}
