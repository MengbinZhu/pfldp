netcdf ropp_testb {
dimensions:
	dim_unlim = UNLIMITED ; // (1 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1a = 1 ;
	dim_lev1b = 293 ;
	dim_lev2a = 273 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 360. ;
	double dtime(dim_unlim, dim_lev1a) ;
		dtime:long_name = "Time since start of occultation" ;
		dtime:units = "seconds" ;
		dtime:valid_range = -1., 240. ;
	float snr_L1ca(dim_unlim, dim_lev1a) ;
		snr_L1ca:long_name = "Signal-to-noise ratio (L1, C/A code)" ;
		snr_L1ca:units = "volt / volt" ;
		snr_L1ca:valid_range = 0., 50000. ;
	float snr_L1p(dim_unlim, dim_lev1a) ;
		snr_L1p:long_name = "Signal-to-noise ratio (L1, P code)" ;
		snr_L1p:units = "volt / volt" ;
		snr_L1p:valid_range = 0., 50000. ;
	float snr_L2p(dim_unlim, dim_lev1a) ;
		snr_L2p:long_name = "Signal-to-noise ratio (L2, P code)" ;
		snr_L2p:units = "volt / volt" ;
		snr_L2p:valid_range = 0., 50000. ;
	double phase_L1(dim_unlim, dim_lev1a) ;
		phase_L1:long_name = "Excess phase (L1)" ;
		phase_L1:units = "metres" ;
		phase_L1:valid_range = -1.e+06, 1.e+06 ;
	double phase_L2(dim_unlim, dim_lev1a) ;
		phase_L2:long_name = "Excess phase (L2)" ;
		phase_L2:units = "metres" ;
		phase_L2:valid_range = -1.e+06, 1.e+06 ;
	double r_gns(dim_unlim, xyz, dim_lev1a) ;
		r_gns:long_name = "GNSS transmitter position" ;
		r_gns:units = "metres" ;
		r_gns:valid_range = -4.3e+07, 4.3e+07 ;
		r_gns:reference_frame = "ECF" ;
	double v_gns(dim_unlim, xyz, dim_lev1a) ;
		v_gns:long_name = "GNSS transmitter velocity" ;
		v_gns:units = "metres / seconds" ;
		v_gns:valid_range = -10000., 10000. ;
		v_gns:reference_frame = "ECI" ;
	double r_leo(dim_unlim, xyz, dim_lev1a) ;
		r_leo:long_name = "LEO transmitter position" ;
		r_leo:units = "metres" ;
		r_leo:valid_range = -1.e+07, 1.e+07 ;
		r_leo:reference_frame = "ECF" ;
	double v_leo(dim_unlim, xyz, dim_lev1a) ;
		v_leo:long_name = "LEO transmitter velocity" ;
		v_leo:units = "metres / seconds" ;
		v_leo:valid_range = -10000., 10000. ;
		v_leo:reference_frame = "ECI" ;
	float phase_qual(dim_unlim, dim_lev1a) ;
		phase_qual:long_name = "Quality value for phase (and SNR)" ;
		phase_qual:units = "percent" ;
		phase_qual:valid_range = 0., 100. ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 360. ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float alt_refrac(dim_unlim, dim_lev2a) ;
		alt_refrac:long_name = "Geometric height above geoid for refractivity" ;
		alt_refrac:units = "metres" ;
		alt_refrac:valid_range = -1000., 1.e+05 ;
	float geop_refrac(dim_unlim, dim_lev2a) ;
		geop_refrac:long_name = "Geopotential height above geoid for refractivity" ;
		geop_refrac:units = "geopotential metres" ;
		geop_refrac:valid_range = -1000., 1.e+05 ;
	double refrac(dim_unlim, dim_lev2a) ;
		refrac:long_name = "Refractivity" ;
		refrac:units = "N-units" ;
		refrac:valid_range = 0., 500. ;
	double refrac_sigma(dim_unlim, dim_lev2a) ;
		refrac_sigma:long_name = "Estimated error (1-sigma) for refractivity" ;
		refrac_sigma:units = "N-units" ;
		refrac_sigma:valid_range = 0., 50. ;
	float refrac_qual(dim_unlim, dim_lev2a) ;
		refrac_qual:long_name = "Quality value for refractivity" ;
		refrac_qual:units = "percent" ;
		refrac_qual:valid_range = 0., 100. ;
	double dry_temp(dim_unlim, dim_lev2a) ;
		dry_temp:long_name = "Dry temperature" ;
		dry_temp:units = "kelvin" ;
		dry_temp:valid_range = 150., 350. ;
	double dry_temp_sigma(dim_unlim, dim_lev2a) ;
		dry_temp_sigma:long_name = "Estimated error (1-sigma) for dry temperature" ;
		dry_temp_sigma:units = "kelvin" ;
		dry_temp_sigma:valid_range = 0., 50. ;
	float dry_temp_qual(dim_unlim, dim_lev2a) ;
		dry_temp_qual:long_name = "Quality value for dry temperature" ;
		dry_temp_qual:units = "percent" ;
		dry_temp_qual:valid_range = 0., 100. ;

// global attributes:
		:title = "ROPP Radio Occultation data" ;
		:institution = "DMI  (ROM SAF)" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "DMI  (ROM SAF)" ;
		:processing_date = "2012-12-12 15:17:20.714" ;
		:pod_method = "UNKNOWN" ;
		:phase_method = "UNKNOWN" ;
		:bangle_method = "UNKNOWN" ;
		:refrac_method = "UNKNOWN" ;
		:meteo_method = "UNKNOWN" ;
		:thin_method = "UNKNOWN" ;
		:software_version = "UNKNOWN" ;
		:_FillValue = -9.9999e+07 ;
data:

 occ_id =
  "OC_20090817215807_META_G027_DMI_" ;

 gns_id =
  "G027" ;

 leo_id =
  "META" ;

 stn_id =
  "UNKN" ;

 start_time = 3.0386e+08 ;

 year = 2009 ;

 month = 8 ;

 day = 17 ;

 hour = 21 ;

 minute = 58 ;

 second = 7 ;

 msec = 814 ;

 pcd = 4 ;

 overall_qual = -9.9999e+07 ;

 time = 3.0386e+08 ;

 time_offset = 5.771 ;

 lat = 50.543 ;

 lon = -3.89 ;

 undulation = 52.5 ;

 roc = 6.3745e+06 ;

 r_coc =
  -3890.3, 9640.6, 20397 ;

 azimuth = -9.9999e+07 ;

 dtime =
  0 ;

 snr_L1ca =
  -9.9999e+07 ;

 snr_L1p =
  -9.9999e+07 ;

 snr_L2p =
  -9.9999e+07 ;

 phase_L1 =
  -9.9999e+07 ;

 phase_L2 =
  -9.9999e+07 ;

 r_gns =
  -9.9999e+07,
  -9.9999e+07,
  -9.9999e+07 ;

 v_gns =
  -9.9999e+07,
  -9.9999e+07,
  -9.9999e+07 ;

 r_leo =
  -9.9999e+07,
  -9.9999e+07,
  -9.9999e+07 ;

 v_leo =
  -9.9999e+07,
  -9.9999e+07,
  -9.9999e+07 ;

 phase_qual =
  -9.9999e+07 ;

 lat_tp =
  50.524, 50.525, 50.527, 50.529, 50.53, 50.532, 50.534, 50.536, 50.538, 
    50.54, 50.542, 50.544, 50.546, 50.547, 50.548, 50.55, 50.551, 50.552, 
    50.554, 50.555, 50.556, 50.558, 50.559, 50.561, 50.562, 50.564, 50.565, 
    50.567, 50.568, 50.57, 50.572, 50.573, 50.574, 50.576, 50.577, 50.578, 
    50.58, 50.581, 50.582, 50.583, 50.584, 50.585, 50.587, 50.588, 50.59, 
    50.591, 50.592, 50.594, 50.595, 50.596, 50.597, 50.598, 50.6, 50.601, 
    50.602, 50.603, 50.605, 50.606, 50.607, 50.608, 50.609, 50.61, 50.611, 
    50.612, 50.613, 50.615, 50.616, 50.617, 50.618, 50.619, 50.62, 50.621, 
    50.622, 50.622, 50.623, 50.624, 50.625, 50.626, 50.627, 50.628, 50.629, 
    50.63, 50.632, 50.633, 50.634, 50.635, 50.636, 50.636, 50.637, 50.638, 
    50.639, 50.64, 50.641, 50.642, 50.643, 50.644, 50.644, 50.645, 50.646, 
    50.647, 50.648, 50.649, 50.65, 50.651, 50.652, 50.653, 50.653, 50.654, 
    50.655, 50.656, 50.657, 50.658, 50.659, 50.66, 50.661, 50.661, 50.662, 
    50.663, 50.664, 50.664, 50.665, 50.666, 50.666, 50.667, 50.668, 50.669, 
    50.67, 50.671, 50.672, 50.673, 50.674, 50.675, 50.676, 50.676, 50.677, 
    50.678, 50.679, 50.68, 50.681, 50.681, 50.682, 50.683, 50.683, 50.684, 
    50.685, 50.686, 50.687, 50.687, 50.688, 50.689, 50.689, 50.69, 50.69, 
    50.691, 50.692, 50.692, 50.694, 50.695, 50.696, 50.697, 50.698, 50.699, 
    50.7, 50.701, 50.701, 50.702, 50.702, 50.703, 50.704, 50.705, 50.706, 
    50.707, 50.707, 50.708, 50.709, 50.71, 50.71, 50.711, 50.711, 50.712, 
    50.713, 50.714, 50.715, 50.716, 50.716, 50.717, 50.718, 50.718, 50.719, 
    50.72, 50.721, 50.722, 50.723, 50.724, 50.725, 50.726, 50.726, 50.727, 
    50.728, 50.728, 50.729, 50.73, 50.731, 50.731, 50.732, 50.733, 50.734, 
    50.734, 50.735, 50.735, 50.736, 50.736, 50.737, 50.738, 50.738, 50.74, 
    50.741, 50.742, 50.743, 50.744, 50.744, 50.745, 50.746, 50.746, 50.747, 
    50.748, 50.748, 50.749, 50.751, 50.752, 50.752, 50.753, 50.754, 50.755, 
    50.755, 50.756, 50.756, 50.757, 50.758, 50.758, 50.759, 50.76, 50.76, 
    50.761, 50.762, 50.763, 50.764, 50.765, 50.766, 50.767, 50.767, 50.768, 
    50.768, 50.769, 50.77, 50.771, 50.772, 50.773, 50.774, 50.774, 50.775, 
    50.775, 50.776, 50.777, 50.778, 50.779, 50.78, 50.78, 50.781, 50.782, 
    50.782, 50.783, 50.784, 50.785, 50.785, 50.786, 50.787, 50.787, 50.788, 
    50.789, 50.79, 50.79, 50.791, 50.792, 50.793, 50.793, 50.794, 50.795, 
    50.796, 50.797, 50.798, 50.799, 50.8 ;

 lon_tp =
  -4.015, -4.018, -4.021, -4.023, -4.026, -4.029, -4.031, -4.034, -4.037, 
    -4.039, -4.042, -4.045, -4.047, -4.05, -4.053, -4.055, -4.058, -4.061, 
    -4.064, -4.066, -4.069, -4.072, -4.075, -4.077, -4.08, -4.083, -4.086, 
    -4.088, -4.091, -4.094, -4.096, -4.099, -4.102, -4.105, -4.107, -4.11, 
    -4.113, -4.116, -4.119, -4.122, -4.124, -4.127, -4.13, -4.133, -4.135, 
    -4.138, -4.141, -4.144, -4.147, -4.149, -4.152, -4.155, -4.158, -4.161, 
    -4.164, -4.166, -4.169, -4.172, -4.175, -4.178, -4.181, -4.184, -4.186, 
    -4.189, -4.192, -4.195, -4.198, -4.201, -4.204, -4.207, -4.21, -4.212, 
    -4.215, -4.218, -4.221, -4.224, -4.227, -4.23, -4.233, -4.236, -4.239, 
    -4.242, -4.244, -4.247, -4.25, -4.253, -4.256, -4.259, -4.262, -4.265, 
    -4.268, -4.271, -4.274, -4.277, -4.28, -4.282, -4.285, -4.288, -4.291, 
    -4.294, -4.297, -4.3, -4.303, -4.306, -4.309, -4.312, -4.315, -4.318, 
    -4.321, -4.324, -4.327, -4.33, -4.333, -4.335, -4.338, -4.341, -4.344, 
    -4.347, -4.35, -4.353, -4.356, -4.359, -4.362, -4.365, -4.368, -4.371, 
    -4.374, -4.377, -4.38, -4.383, -4.386, -4.389, -4.392, -4.395, -4.398, 
    -4.401, -4.404, -4.406, -4.409, -4.412, -4.415, -4.418, -4.421, -4.424, 
    -4.427, -4.43, -4.433, -4.436, -4.439, -4.442, -4.445, -4.448, -4.451, 
    -4.454, -4.457, -4.46, -4.463, -4.466, -4.469, -4.472, -4.475, -4.478, 
    -4.481, -4.484, -4.487, -4.49, -4.493, -4.496, -4.499, -4.502, -4.504, 
    -4.507, -4.51, -4.513, -4.516, -4.519, -4.522, -4.525, -4.528, -4.531, 
    -4.534, -4.537, -4.54, -4.543, -4.546, -4.549, -4.552, -4.555, -4.558, 
    -4.561, -4.564, -4.567, -4.57, -4.573, -4.576, -4.579, -4.582, -4.585, 
    -4.588, -4.591, -4.594, -4.596, -4.599, -4.602, -4.605, -4.608, -4.611, 
    -4.614, -4.617, -4.62, -4.623, -4.626, -4.629, -4.632, -4.635, -4.638, 
    -4.641, -4.644, -4.647, -4.65, -4.653, -4.656, -4.659, -4.662, -4.665, 
    -4.668, -4.671, -4.674, -4.677, -4.679, -4.682, -4.685, -4.688, -4.691, 
    -4.694, -4.697, -4.7, -4.703, -4.706, -4.709, -4.712, -4.715, -4.718, 
    -4.721, -4.724, -4.727, -4.73, -4.733, -4.736, -4.739, -4.742, -4.745, 
    -4.748, -4.751, -4.754, -4.757, -4.76, -4.762, -4.765, -4.768, -4.771, 
    -4.774, -4.777, -4.78, -4.783, -4.786, -4.789, -4.792, -4.795, -4.798, 
    -4.801, -4.804, -4.807, -4.81, -4.813, -4.816, -4.819, -4.822, -4.825, 
    -4.828, -4.831, -4.834, -4.836, -4.839, -4.842, -4.845, -4.848, -4.851, 
    -4.854, -4.857, -4.86, -4.863, -4.866 ;

 azimuth_tp =
  193.13, 193.13, 193.13, 193.13, 193.12, 193.12, 193.12, 193.12, 193.12, 
    193.12, 193.11, 193.11, 193.11, 193.11, 193.1, 193.1, 193.1, 193.1, 
    193.1, 193.09, 193.09, 193.09, 193.09, 193.09, 193.08, 193.08, 193.08, 
    193.08, 193.08, 193.07, 193.07, 193.07, 193.07, 193.07, 193.06, 193.06, 
    193.06, 193.06, 193.05, 193.05, 193.05, 193.05, 193.05, 193.04, 193.04, 
    193.04, 193.04, 193.04, 193.03, 193.03, 193.03, 193.03, 193.03, 193.02, 
    193.02, 193.02, 193.02, 193.01, 193.01, 193.01, 193.01, 193.01, 193, 193, 
    193, 193, 193, 192.99, 192.99, 192.99, 192.99, 192.98, 192.98, 192.98, 
    192.98, 192.98, 192.97, 192.97, 192.97, 192.97, 192.96, 192.96, 192.96, 
    192.96, 192.96, 192.95, 192.95, 192.95, 192.95, 192.94, 192.94, 192.94, 
    192.94, 192.94, 192.93, 192.93, 192.93, 192.93, 192.92, 192.92, 192.92, 
    192.92, 192.92, 192.91, 192.91, 192.91, 192.91, 192.9, 192.9, 192.9, 
    192.9, 192.9, 192.89, 192.89, 192.89, 192.89, 192.88, 192.88, 192.88, 
    192.88, 192.88, 192.87, 192.87, 192.87, 192.87, 192.86, 192.86, 192.86, 
    192.86, 192.86, 192.85, 192.85, 192.85, 192.85, 192.84, 192.84, 192.84, 
    192.84, 192.84, 192.83, 192.83, 192.83, 192.83, 192.82, 192.82, 192.82, 
    192.82, 192.81, 192.81, 192.81, 192.81, 192.81, 192.8, 192.8, 192.8, 
    192.8, 192.79, 192.79, 192.79, 192.79, 192.79, 192.78, 192.78, 192.78, 
    192.78, 192.77, 192.77, 192.77, 192.77, 192.76, 192.76, 192.76, 192.76, 
    192.76, 192.75, 192.75, 192.75, 192.75, 192.75, 192.74, 192.74, 192.74, 
    192.74, 192.73, 192.73, 192.73, 192.73, 192.72, 192.72, 192.72, 192.72, 
    192.72, 192.71, 192.71, 192.71, 192.71, 192.7, 192.7, 192.7, 192.7, 
    192.7, 192.69, 192.69, 192.69, 192.69, 192.68, 192.68, 192.68, 192.68, 
    192.68, 192.67, 192.67, 192.67, 192.67, 192.66, 192.66, 192.66, 192.66, 
    192.65, 192.65, 192.65, 192.65, 192.65, 192.64, 192.64, 192.64, 192.64, 
    192.63, 192.63, 192.63, 192.63, 192.63, 192.62, 192.62, 192.62, 192.62, 
    192.61, 192.61, 192.61, 192.61, 192.61, 192.6, 192.6, 192.6, 192.6, 
    192.59, 192.59, 192.59, 192.59, 192.59, 192.58, 192.58, 192.58, 192.58, 
    192.57, 192.57, 192.57, 192.57, 192.57, 192.56, 192.56, 192.56, 192.56, 
    192.55, 192.55, 192.55, 192.55, 192.54, 192.54, 192.54, 192.54, 192.54, 
    192.53, 192.53, 192.53, 192.53, 192.52, 192.52, 192.52, 192.52, 192.52, 
    192.51, 192.51, 192.51, 192.51, 192.5, 192.5, 192.5, 192.5, 192.5, 
    192.49, 192.49, 192.49 ;

 impact_L1 =
  6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3768e+06, 6.3768e+06, 
    6.377e+06, 6.3773e+06, 6.3776e+06, 6.3778e+06, 6.3779e+06, 6.3779e+06, 
    6.378e+06, 6.378e+06, 6.3781e+06, 6.3783e+06, 6.3786e+06, 6.3788e+06, 
    6.379e+06, 6.379e+06, 6.3788e+06, 6.3786e+06, 6.3785e+06, 6.3784e+06, 
    6.3782e+06, 6.3781e+06, 6.378e+06, 6.3781e+06, 6.3784e+06, 6.3788e+06, 
    6.3791e+06, 6.3793e+06, 6.3793e+06, 6.3792e+06, 6.379e+06, 6.3789e+06, 
    6.3787e+06, 6.3787e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3789e+06, 
    6.3791e+06, 6.3793e+06, 6.3792e+06, 6.3791e+06, 6.3789e+06, 6.3788e+06, 
    6.379e+06, 6.3793e+06, 6.3794e+06, 6.3793e+06, 6.3793e+06, 6.3791e+06, 
    6.379e+06, 6.3791e+06, 6.3793e+06, 6.3795e+06, 6.3798e+06, 6.38e+06, 
    6.38e+06, 6.3798e+06, 6.3795e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3805e+06, 6.3807e+06, 6.381e+06, 6.3811e+06, 
    6.3812e+06, 6.3812e+06, 6.3813e+06, 6.3814e+06, 6.3815e+06, 6.3816e+06, 
    6.3817e+06, 6.3819e+06, 6.382e+06, 6.3821e+06, 6.3822e+06, 6.3823e+06, 
    6.3824e+06, 6.3825e+06, 6.3826e+06, 6.3827e+06, 6.3829e+06, 6.383e+06, 
    6.3831e+06, 6.3833e+06, 6.3833e+06, 6.3834e+06, 6.3835e+06, 6.3836e+06, 
    6.3837e+06, 6.3838e+06, 6.3839e+06, 6.3841e+06, 6.3842e+06, 6.3844e+06, 
    6.3846e+06, 6.3848e+06, 6.3849e+06, 6.385e+06, 6.3851e+06, 6.3852e+06, 
    6.3854e+06, 6.3855e+06, 6.3856e+06, 6.3858e+06, 6.3859e+06, 6.3861e+06, 
    6.3863e+06, 6.3864e+06, 6.3865e+06, 6.3867e+06, 6.387e+06, 6.3872e+06, 
    6.3875e+06, 6.3876e+06, 6.3878e+06, 6.3879e+06, 6.388e+06, 6.3881e+06, 
    6.3882e+06, 6.3883e+06, 6.3884e+06, 6.3885e+06, 6.3886e+06, 6.3887e+06, 
    6.3887e+06, 6.3888e+06, 6.389e+06, 6.3891e+06, 6.3892e+06, 6.3893e+06, 
    6.3894e+06, 6.3895e+06, 6.3897e+06, 6.3899e+06, 6.39e+06, 6.3902e+06, 
    6.3903e+06, 6.3904e+06, 6.3906e+06, 6.3908e+06, 6.3909e+06, 6.391e+06, 
    6.3912e+06, 6.3914e+06, 6.3916e+06, 6.3918e+06, 6.392e+06, 6.3922e+06, 
    6.3923e+06, 6.3925e+06, 6.3927e+06, 6.3929e+06, 6.3931e+06, 6.3933e+06, 
    6.3935e+06, 6.3937e+06, 6.3939e+06, 6.3941e+06, 6.3943e+06, 6.3945e+06, 
    6.3948e+06, 6.395e+06, 6.3953e+06, 6.3955e+06, 6.3958e+06, 6.396e+06, 
    6.3963e+06, 6.3966e+06, 6.3968e+06, 6.3971e+06, 6.3973e+06, 6.3976e+06, 
    6.3979e+06, 6.3982e+06, 6.3985e+06, 6.3988e+06, 6.3991e+06, 6.3994e+06, 
    6.3997e+06, 6.4e+06, 6.4003e+06, 6.4006e+06, 6.4009e+06, 6.4013e+06, 
    6.4016e+06, 6.4019e+06, 6.4022e+06, 6.4026e+06, 6.403e+06, 6.4033e+06, 
    6.4036e+06, 6.404e+06, 6.4044e+06, 6.4047e+06, 6.4051e+06, 6.4055e+06, 
    6.4058e+06, 6.4062e+06, 6.4066e+06, 6.4069e+06, 6.4073e+06, 6.4076e+06, 
    6.408e+06, 6.4084e+06, 6.4088e+06, 6.4092e+06, 6.4096e+06, 6.41e+06, 
    6.4104e+06, 6.4108e+06, 6.4111e+06, 6.4115e+06, 6.4119e+06, 6.4123e+06, 
    6.4127e+06, 6.4131e+06, 6.4135e+06, 6.4139e+06, 6.4143e+06, 6.4147e+06, 
    6.4151e+06, 6.4155e+06, 6.4159e+06, 6.4163e+06, 6.4167e+06, 6.4171e+06, 
    6.4175e+06, 6.4179e+06, 6.4183e+06, 6.4187e+06, 6.4191e+06, 6.4195e+06, 
    6.4199e+06, 6.4203e+06, 6.4207e+06, 6.4211e+06, 6.4215e+06, 6.4219e+06, 
    6.4224e+06, 6.4228e+06, 6.4232e+06, 6.4236e+06, 6.424e+06, 6.4243e+06, 
    6.4247e+06, 6.4252e+06, 6.4256e+06, 6.426e+06, 6.4264e+06, 6.4268e+06, 
    6.4272e+06, 6.4276e+06, 6.428e+06, 6.4284e+06, 6.4289e+06, 6.4293e+06, 
    6.4297e+06, 6.4301e+06, 6.4305e+06, 6.4309e+06, 6.4313e+06, 6.4317e+06, 
    6.4321e+06, 6.4325e+06, 6.4329e+06, 6.4333e+06, 6.4337e+06, 6.4341e+06, 
    6.4345e+06, 6.4349e+06, 6.4354e+06, 6.4358e+06, 6.4362e+06, 6.4367e+06, 
    6.4371e+06, 6.4374e+06, 6.4378e+06, 6.4382e+06, 6.4386e+06, 6.439e+06, 
    6.4395e+06, 6.4399e+06, 6.4402e+06, 6.4406e+06, 6.441e+06 ;

 impact_L2 =
  6.3923e+06, 6.3923e+06, 6.3924e+06, 6.3926e+06, 6.3927e+06, 6.3928e+06, 
    6.3929e+06, 6.393e+06, 6.3931e+06, 6.3932e+06, 6.3934e+06, 6.3935e+06, 
    6.3936e+06, 6.3937e+06, 6.3938e+06, 6.3939e+06, 6.394e+06, 6.3941e+06, 
    6.3942e+06, 6.3943e+06, 6.3944e+06, 6.3946e+06, 6.3947e+06, 6.3949e+06, 
    6.3951e+06, 6.3952e+06, 6.3954e+06, 6.3955e+06, 6.3957e+06, 6.3958e+06, 
    6.396e+06, 6.3961e+06, 6.3963e+06, 6.3964e+06, 6.3965e+06, 6.3967e+06, 
    6.3968e+06, 6.397e+06, 6.3971e+06, 6.3973e+06, 6.3974e+06, 6.3976e+06, 
    6.3977e+06, 6.3979e+06, 6.3981e+06, 6.3983e+06, 6.3985e+06, 6.3987e+06, 
    6.3988e+06, 6.399e+06, 6.3992e+06, 6.3993e+06, 6.3995e+06, 6.3996e+06, 
    6.3998e+06, 6.3999e+06, 6.4001e+06, 6.4003e+06, 6.4005e+06, 6.4007e+06, 
    6.4009e+06, 6.4011e+06, 6.4012e+06, 6.4014e+06, 6.4016e+06, 6.4018e+06, 
    6.402e+06, 6.4022e+06, 6.4024e+06, 6.4026e+06, 6.4028e+06, 6.403e+06, 
    6.4032e+06, 6.4034e+06, 6.4036e+06, 6.4038e+06, 6.404e+06, 6.4042e+06, 
    6.4044e+06, 6.4046e+06, 6.4048e+06, 6.405e+06, 6.4052e+06, 6.4055e+06, 
    6.4057e+06, 6.4059e+06, 6.4061e+06, 6.4063e+06, 6.4065e+06, 6.4067e+06, 
    6.4069e+06, 6.4071e+06, 6.4073e+06, 6.4075e+06, 6.4077e+06, 6.408e+06, 
    6.4082e+06, 6.4084e+06, 6.4086e+06, 6.4088e+06, 6.4091e+06, 6.4093e+06, 
    6.4095e+06, 6.4097e+06, 6.41e+06, 6.4102e+06, 6.4104e+06, 6.4106e+06, 
    6.4108e+06, 6.4111e+06, 6.4113e+06, 6.4115e+06, 6.4117e+06, 6.4119e+06, 
    6.4122e+06, 6.4124e+06, 6.4126e+06, 6.4128e+06, 6.4131e+06, 6.4133e+06, 
    6.4135e+06, 6.4137e+06, 6.4139e+06, 6.4142e+06, 6.4144e+06, 6.4146e+06, 
    6.4149e+06, 6.4151e+06, 6.4154e+06, 6.4156e+06, 6.4158e+06, 6.4161e+06, 
    6.4163e+06, 6.4165e+06, 6.4167e+06, 6.4169e+06, 6.4172e+06, 6.4174e+06, 
    6.4176e+06, 6.4178e+06, 6.4181e+06, 6.4183e+06, 6.4185e+06, 6.4187e+06, 
    6.419e+06, 6.4192e+06, 6.4194e+06, 6.4197e+06, 6.4199e+06, 6.4202e+06, 
    6.4204e+06, 6.4206e+06, 6.4209e+06, 6.4211e+06, 6.4213e+06, 6.4216e+06, 
    6.4218e+06, 6.422e+06, 6.4223e+06, 6.4226e+06, 6.4228e+06, 6.4231e+06, 
    6.4233e+06, 6.4235e+06, 6.4237e+06, 6.4239e+06, 6.4241e+06, 6.4243e+06, 
    6.4245e+06, 6.4247e+06, 6.425e+06, 6.4252e+06, 6.4255e+06, 6.4257e+06, 
    6.426e+06, 6.4262e+06, 6.4264e+06, 6.4267e+06, 6.4269e+06, 6.4271e+06, 
    6.4273e+06, 6.4276e+06, 6.4278e+06, 6.428e+06, 6.4283e+06, 6.4285e+06, 
    6.4288e+06, 6.429e+06, 6.4293e+06, 6.4295e+06, 6.4297e+06, 6.4299e+06, 
    6.4302e+06, 6.4304e+06, 6.4307e+06, 6.4309e+06, 6.4311e+06, 6.4314e+06, 
    6.4316e+06, 6.4318e+06, 6.432e+06, 6.4322e+06, 6.4324e+06, 6.4327e+06, 
    6.4329e+06, 6.4332e+06, 6.4334e+06, 6.4336e+06, 6.4339e+06, 6.4341e+06, 
    6.4343e+06, 6.4346e+06, 6.4348e+06, 6.435e+06, 6.4353e+06, 6.4355e+06, 
    6.4358e+06, 6.436e+06, 6.4363e+06, 6.4366e+06, 6.4368e+06, 6.437e+06, 
    6.4372e+06, 6.4374e+06, 6.4376e+06, 6.4379e+06, 6.4381e+06, 6.4383e+06, 
    6.4385e+06, 6.4388e+06, 6.439e+06, 6.4393e+06, 6.4395e+06, 6.4397e+06, 
    6.44e+06, 6.4402e+06, 6.4404e+06, 6.4406e+06, 6.4408e+06, 6.441e+06, 
    6.4413e+06, 6.4415e+06, 6.4418e+06, 6.442e+06, 6.4423e+06, 6.4425e+06, 
    6.4428e+06, 6.443e+06, 6.4432e+06, 6.4435e+06, 6.4437e+06, 6.4439e+06, 
    6.4441e+06, 6.4443e+06, 6.4445e+06, 6.4448e+06, 6.445e+06, 6.4453e+06, 
    6.4455e+06, 6.4458e+06, 6.446e+06, 6.4462e+06, 6.4464e+06, 6.4466e+06, 
    6.4469e+06, 6.4471e+06, 6.4473e+06, 6.4476e+06, 6.4478e+06, 6.4481e+06, 
    6.4483e+06, 6.4485e+06, 6.4487e+06, 6.449e+06, 6.4492e+06, 6.4494e+06, 
    6.4497e+06, 6.4499e+06, 6.4501e+06, 6.4504e+06, 6.4506e+06, 6.4508e+06, 
    6.4511e+06, 6.4513e+06, 6.4515e+06, 6.4518e+06, 6.452e+06, 6.4522e+06, 
    6.4525e+06, 6.4527e+06, 6.4529e+06, 6.4531e+06, 6.4534e+06 ;

 impact =
  6.393e+06, 6.3931e+06, 6.3933e+06, 6.3934e+06, 6.3935e+06, 6.3936e+06, 
    6.3937e+06, 6.3939e+06, 6.394e+06, 6.3941e+06, 6.3942e+06, 6.3943e+06, 
    6.3944e+06, 6.3945e+06, 6.3947e+06, 6.3948e+06, 6.395e+06, 6.3951e+06, 
    6.3953e+06, 6.3954e+06, 6.3956e+06, 6.3957e+06, 6.3959e+06, 6.396e+06, 
    6.3961e+06, 6.3963e+06, 6.3964e+06, 6.3966e+06, 6.3967e+06, 6.3969e+06, 
    6.397e+06, 6.3972e+06, 6.3973e+06, 6.3975e+06, 6.3976e+06, 6.3978e+06, 
    6.398e+06, 6.3982e+06, 6.3984e+06, 6.3985e+06, 6.3987e+06, 6.3989e+06, 
    6.399e+06, 6.3992e+06, 6.3994e+06, 6.3995e+06, 6.3997e+06, 6.3998e+06, 
    6.4e+06, 6.4002e+06, 6.4004e+06, 6.4006e+06, 6.4008e+06, 6.4009e+06, 
    6.4011e+06, 6.4013e+06, 6.4015e+06, 6.4017e+06, 6.4019e+06, 6.4021e+06, 
    6.4022e+06, 6.4025e+06, 6.4027e+06, 6.4029e+06, 6.403e+06, 6.4032e+06, 
    6.4034e+06, 6.4036e+06, 6.4038e+06, 6.404e+06, 6.4042e+06, 6.4045e+06, 
    6.4047e+06, 6.4049e+06, 6.4051e+06, 6.4053e+06, 6.4055e+06, 6.4057e+06, 
    6.406e+06, 6.4062e+06, 6.4064e+06, 6.4066e+06, 6.4068e+06, 6.407e+06, 
    6.4072e+06, 6.4074e+06, 6.4076e+06, 6.4078e+06, 6.408e+06, 6.4083e+06, 
    6.4085e+06, 6.4087e+06, 6.4089e+06, 6.4091e+06, 6.4094e+06, 6.4096e+06, 
    6.4098e+06, 6.41e+06, 6.4103e+06, 6.4105e+06, 6.4107e+06, 6.4109e+06, 
    6.4111e+06, 6.4114e+06, 6.4116e+06, 6.4118e+06, 6.412e+06, 6.4123e+06, 
    6.4125e+06, 6.4127e+06, 6.4129e+06, 6.4132e+06, 6.4134e+06, 6.4136e+06, 
    6.4138e+06, 6.414e+06, 6.4143e+06, 6.4145e+06, 6.4147e+06, 6.415e+06, 
    6.4152e+06, 6.4154e+06, 6.4157e+06, 6.4159e+06, 6.4161e+06, 6.4164e+06, 
    6.4166e+06, 6.4168e+06, 6.417e+06, 6.4172e+06, 6.4175e+06, 6.4177e+06, 
    6.4179e+06, 6.4182e+06, 6.4184e+06, 6.4186e+06, 6.4188e+06, 6.4191e+06, 
    6.4193e+06, 6.4195e+06, 6.4198e+06, 6.42e+06, 6.4202e+06, 6.4205e+06, 
    6.4207e+06, 6.421e+06, 6.4212e+06, 6.4214e+06, 6.4216e+06, 6.4219e+06, 
    6.4221e+06, 6.4224e+06, 6.4226e+06, 6.4229e+06, 6.4231e+06, 6.4233e+06, 
    6.4236e+06, 6.4238e+06, 6.424e+06, 6.4242e+06, 6.4244e+06, 6.4246e+06, 
    6.4249e+06, 6.4251e+06, 6.4254e+06, 6.4256e+06, 6.4258e+06, 6.4261e+06, 
    6.4263e+06, 6.4265e+06, 6.4268e+06, 6.427e+06, 6.4272e+06, 6.4274e+06, 
    6.4277e+06, 6.4279e+06, 6.4281e+06, 6.4284e+06, 6.4286e+06, 6.4289e+06, 
    6.4291e+06, 6.4293e+06, 6.4296e+06, 6.4298e+06, 6.43e+06, 6.4303e+06, 
    6.4305e+06, 6.4307e+06, 6.431e+06, 6.4312e+06, 6.4314e+06, 6.4317e+06, 
    6.4319e+06, 6.4321e+06, 6.4323e+06, 6.4326e+06, 6.4328e+06, 6.433e+06, 
    6.4333e+06, 6.4335e+06, 6.4337e+06, 6.434e+06, 6.4342e+06, 6.4344e+06, 
    6.4347e+06, 6.4349e+06, 6.4351e+06, 6.4354e+06, 6.4356e+06, 6.4359e+06, 
    6.4361e+06, 6.4364e+06, 6.4366e+06, 6.4368e+06, 6.4371e+06, 6.4373e+06, 
    6.4375e+06, 6.4377e+06, 6.4379e+06, 6.4382e+06, 6.4384e+06, 6.4386e+06, 
    6.4389e+06, 6.4391e+06, 6.4393e+06, 6.4396e+06, 6.4398e+06, 6.44e+06, 
    6.4402e+06, 6.4405e+06, 6.4407e+06, 6.4409e+06, 6.4411e+06, 6.4414e+06, 
    6.4416e+06, 6.4419e+06, 6.4421e+06, 6.4423e+06, 6.4426e+06, 6.4428e+06, 
    6.4431e+06, 6.4433e+06, 6.4435e+06, 6.4438e+06, 6.444e+06, 6.4442e+06, 
    6.4444e+06, 6.4446e+06, 6.4449e+06, 6.4451e+06, 6.4453e+06, 6.4456e+06, 
    6.4458e+06, 6.4461e+06, 6.4463e+06, 6.4465e+06, 6.4467e+06, 6.447e+06, 
    6.4472e+06, 6.4474e+06, 6.4477e+06, 6.4479e+06, 6.4481e+06, 6.4484e+06, 
    6.4486e+06, 6.4488e+06, 6.449e+06, 6.4493e+06, 6.4495e+06, 6.4497e+06, 
    6.45e+06, 6.4502e+06, 6.4504e+06, 6.4507e+06, 6.4509e+06, 6.4511e+06, 
    6.4514e+06, 6.4516e+06, 6.4518e+06, 6.4521e+06, 6.4523e+06, 6.4525e+06, 
    6.4527e+06, 6.453e+06, 6.4532e+06, 6.4535e+06, 6.4537e+06, 6.4539e+06, 
    6.4541e+06, 6.4544e+06, 6.4546e+06, 6.4548e+06, 6.455e+06 ;

 impact_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1 =
  0.022189, 0.022057, 0.021921, 0.021764, 0.021609, 0.021478, 0.021393, 
    0.021346, 0.021305, 0.021237, 0.021124, 0.021, 0.020882, 0.020749, 
    0.020636, 0.020557, 0.02051, 0.020461, 0.02037, 0.020235, 0.020031, 
    0.019822, 0.019623, 0.019447, 0.019257, 0.019065, 0.018903, 0.018783, 
    0.018748, 0.018742, 0.018711, 0.018626, 0.018501, 0.018327, 0.018119, 
    0.017923, 0.017735, 0.017576, 0.017478, 0.017335, 0.01719, 0.017088, 
    0.017012, 0.016928, 0.016761, 0.016583, 0.016375, 0.016215, 0.016146, 
    0.016081, 0.015977, 0.015826, 0.015659, 0.015461, 0.015301, 0.015188, 
    0.015096, 0.015029, 0.014987, 0.014903, 0.014765, 0.014565, 0.014325, 
    0.011613, 0.011476, 0.011328, 0.011165, 0.011031, 0.010936, 0.010864, 
    0.010805, 0.010719, 0.010604, 0.010474, 0.01036, 0.010242, 0.010133, 
    0.010035, 0.0099327, 0.0098332, 0.0097326, 0.009623, 0.0095129, 
    0.0094044, 0.0093058, 0.0091953, 0.009089, 0.0089935, 0.0089037, 
    0.0088037, 0.0087075, 0.008614, 0.0085003, 0.0083881, 0.0082711, 
    0.0081527, 0.0080389, 0.0079446, 0.0078476, 0.0077479, 0.0076585, 
    0.0075791, 0.0075031, 0.0074206, 0.0073261, 0.0072201, 0.0071161, 
    0.0070176, 0.0069219, 0.0068267, 0.006732, 0.0066394, 0.0065526, 
    0.0064699, 0.0063798, 0.0062847, 0.00619, 0.0061141, 0.0060544, 
    0.0059994, 0.0059347, 0.0058525, 0.0057552, 0.0056494, 0.0055458, 
    0.0054368, 0.0053254, 0.0052184, 0.0051143, 0.0050071, 0.0048978, 
    0.0047818, 0.0046666, 0.0045633, 0.0044714, 0.0043756, 0.0042704, 
    0.0041611, 0.0040499, 0.0039527, 0.0038642, 0.0037761, 0.0036845, 
    0.003593, 0.0035012, 0.0034108, 0.0033233, 0.0032311, 0.0031386, 
    0.0030475, 0.0029568, 0.0028731, 0.0027984, 0.0027258, 0.0026527, 
    0.002578, 0.0024982, 0.0024178, 0.002338, 0.0022585, 0.0021828, 
    0.0021143, 0.0020465, 0.0019766, 0.0019013, 0.0018215, 0.0017448, 
    0.0016775, 0.0016211, 0.0015672, 0.0015134, 0.0014584, 0.0014033, 
    0.0013501, 0.0012979, 0.0012456, 0.0011909, 0.0011363, 0.0010832, 
    0.0010358, 0.00099604, 0.00096376, 0.00093145, 0.00089331, 0.00084703, 
    0.0007971, 0.00074887, 0.00070698, 0.00067412, 0.00064593, 0.00061649, 
    0.00058277, 0.00055106, 0.00052189, 0.00049789, 0.00047699, 0.00045473, 
    0.00042914, 0.00040504, 0.00038479, 0.00036749, 0.00035265, 0.00033951, 
    0.00032677, 0.00031401, 0.00029698, 0.00027567, 0.00025368, 0.00023507, 
    0.00022266, 0.00021463, 0.00020775, 0.00019745, 0.00018616, 0.00017687, 
    0.00017052, 0.00016488, 0.00015671, 0.00014618, 0.00013601, 0.0001284, 
    0.0001231, 0.00011817, 0.00011042, 0.00010135, 9.38e-05, 8.729e-05, 
    8.431e-05, 8.614e-05, 8.908e-05, 8.793e-05, 8.364e-05, 7.558e-05, 
    6.589e-05, 5.871e-05, 5.451e-05, 5.102e-05, 4.686e-05, 4.471e-05, 
    4.47e-05, 4.504e-05, 4.547e-05, 4.615e-05, 4.556e-05, 4.214e-05, 
    4.204e-05, 5.02e-05, 6.025e-05, 6.279e-05, 5.529e-05, 3.961e-05, 
    2.474e-05, 2.094e-05, 2.54e-05, 3.17e-05, 3.512e-05, 3.333e-05, 
    2.727e-05, 2.336e-05, 2.191e-05, 2.262e-05, 2.908e-05, 3.637e-05, 
    3.456e-05, 2.984e-05, 2.807e-05, 3.07e-05, 3.341e-05, 3.476e-05, 
    3.05e-05, 2.114e-05, 1.502e-05, 1.517e-05, 2.015e-05, 2.103e-05, 
    2.12e-05, 1.812e-05, 1.796e-05, 2.145e-05, 3.011e-05, 3.991e-05, 
    4.688e-05, 4.609e-05, 3.367e-05, 2.439e-05, 2.047e-05, 1.985e-05, 
    2.603e-05, 3.228e-05, 2.997e-05, 1.92e-05, 1.222e-05, 1.066e-05 ;

 bangle_L2 =
  0.002548, 0.0025006, 0.0024541, 0.0024094, 0.0023646, 0.0023201, 0.0022776, 
    0.0022348, 0.0021955, 0.0021598, 0.0021231, 0.002085, 0.0020446, 
    0.0020016, 0.0019546, 0.0019047, 0.0018521, 0.0017996, 0.001751, 
    0.0017082, 0.0016722, 0.0016415, 0.0016142, 0.0015879, 0.0015617, 
    0.0015341, 0.001505, 0.0014751, 0.0014452, 0.0014151, 0.0013846, 
    0.0013537, 0.0013222, 0.0012901, 0.0012568, 0.0012239, 0.0011914, 
    0.0011589, 0.0011279, 0.0010986, 0.0010706, 0.0010447, 0.0010209, 
    0.00099968, 0.00098165, 0.00096496, 0.00094779, 0.00092929, 0.00090893, 
    0.00088509, 0.00085803, 0.00082974, 0.00080024, 0.00077059, 0.00074344, 
    0.00071978, 0.0006995, 0.0006829, 0.00066822, 0.00065331, 0.00063712, 
    0.00061757, 0.00059629, 0.00057507, 0.00055557, 0.00053717, 0.00052065, 
    0.00050712, 0.00049618, 0.00048562, 0.00047399, 0.00046141, 0.00044647, 
    0.00043144, 0.00041787, 0.00040545, 0.00039429, 0.00038523, 0.00037665, 
    0.00036803, 0.00036162, 0.00035662, 0.000351, 0.00034491, 0.00033873, 
    0.0003317, 0.00032182, 0.00030986, 0.00029527, 0.00027992, 0.0002658, 
    0.00025222, 0.00024123, 0.00023435, 0.00022962, 0.00022579, 0.00022288, 
    0.00022036, 0.00021562, 0.00020896, 0.00020196, 0.00019512, 0.00018973, 
    0.0001862, 0.00018335, 0.000181, 0.00017841, 0.00017452, 0.00016777, 
    0.00016058, 0.00015359, 0.00014673, 0.00014139, 0.00013763, 0.00013516, 
    0.00013325, 0.00013088, 0.0001275, 0.00012233, 0.00011578, 0.00010966, 
    0.00010405, 9.929e-05, 9.535e-05, 9.282e-05, 9.243e-05, 9.492e-05, 
    9.911e-05, 0.00010375, 0.00010587, 0.00010625, 0.00010426, 0.00010131, 
    9.588e-05, 8.895e-05, 8.054e-05, 7.343e-05, 6.758e-05, 6.366e-05, 
    6.108e-05, 5.86e-05, 5.572e-05, 5.256e-05, 5.012e-05, 4.944e-05, 
    4.963e-05, 5e-05, 5.089e-05, 5.222e-05, 5.328e-05, 5.51e-05, 5.596e-05, 
    5.697e-05, 5.611e-05, 5.339e-05, 5.139e-05, 5.208e-05, 5.56e-05, 
    6.288e-05, 7.292e-05, 8.298e-05, 8.944e-05, 8.961e-05, 8.376e-05, 
    7.224e-05, 5.802e-05, 4.265e-05, 3.038e-05, 2.364e-05, 2.224e-05, 
    2.475e-05, 3.106e-05, 3.865e-05, 4.407e-05, 4.701e-05, 4.69e-05, 
    4.455e-05, 3.99e-05, 3.479e-05, 3.103e-05, 2.827e-05, 2.695e-05, 
    2.69e-05, 2.94e-05, 3.48e-05, 4.273e-05, 5.045e-05, 5.285e-05, 5.063e-05, 
    4.637e-05, 4.199e-05, 3.954e-05, 4.081e-05, 4.393e-05, 4.733e-05, 
    4.996e-05, 5.194e-05, 5.131e-05, 4.835e-05, 4.245e-05, 3.196e-05, 
    2.322e-05, 1.95e-05, 1.845e-05, 2.037e-05, 2.493e-05, 2.894e-05, 
    3.047e-05, 3.149e-05, 3.042e-05, 2.792e-05, 2.647e-05, 2.716e-05, 
    2.757e-05, 2.996e-05, 3.644e-05, 4.556e-05, 5.544e-05, 6.471e-05, 
    7.185e-05, 7.512e-05, 7.433e-05, 6.693e-05, 5.479e-05, 4.427e-05, 
    3.771e-05, 3.197e-05, 2.791e-05, 2.981e-05, 3.422e-05, 4.041e-05, 
    4.554e-05, 4.947e-05, 4.952e-05, 4.393e-05, 3.441e-05, 2.482e-05, 
    1.831e-05, 1.643e-05, 1.398e-05, 1.705e-05, 2.492e-05, 3.187e-05, 
    3.646e-05, 3.983e-05, 4.39e-05, 4.982e-05, 5.43e-05, 5.752e-05, 
    5.948e-05, 5.888e-05, 5.442e-05, 4.431e-05, 3.3e-05, 2.486e-05, 
    2.078e-05, 2.378e-05, 3.149e-05, 4.12e-05, 4.807e-05, 4.779e-05, 
    4.373e-05, 3.762e-05, 3.159e-05, 2.721e-05, 2.65e-05, 2.951e-05, 
    3.409e-05, 3.684e-05, 3.778e-05, 3.605e-05, 3.322e-05, 3.015e-05, 
    2.812e-05, 2.951e-05, 3.319e-05, 3.547e-05, 3.736e-05, 3.782e-05, 
    3.738e-05, 3.681e-05, 3.695e-05, 3.912e-05, 4.28e-05, 4.649e-05, 
    5.128e-05, 5.166e-05, 4.871e-05, 4.46e-05, 4.065e-05, 3.899e-05, 
    4.238e-05, 4.936e-05 ;

 bangle =
  0.0021696, 0.0021214, 0.0020741, 0.0020307, 0.0019901, 0.0019529, 
    0.0019218, 0.0018967, 0.0018789, 0.0018637, 0.0018348, 0.0017945, 
    0.001748, 0.0017016, 0.0016574, 0.0016156, 0.0015754, 0.0015363, 
    0.0014986, 0.0014621, 0.0014258, 0.0013912, 0.0013586, 0.0013292, 
    0.0013019, 0.001277, 0.0012539, 0.0012307, 0.0012042, 0.0011759, 
    0.0011452, 0.001113, 0.0010806, 0.001051, 0.0010241, 0.00099995, 
    0.00097859, 0.0009582, 0.00093786, 0.00091593, 0.0008916, 0.00086437, 
    0.00083595, 0.00080699, 0.00077893, 0.00075371, 0.00073031, 0.00070805, 
    0.00068692, 0.00066691, 0.00064737, 0.0006287, 0.00061077, 0.0005938, 
    0.00057777, 0.00056301, 0.000549, 0.00053468, 0.00052042, 0.0005061, 
    0.00049175, 0.00047758, 0.00046319, 0.00044912, 0.0004351, 0.00042115, 
    0.00040723, 0.00039372, 0.0003812, 0.00036926, 0.0003579, 0.00034721, 
    0.00033674, 0.00032637, 0.00031628, 0.00030661, 0.00029722, 0.00028794, 
    0.00027874, 0.00026995, 0.00026132, 0.00025301, 0.00024448, 0.00023591, 
    0.00022778, 0.00021966, 0.00021208, 0.00020522, 0.00019896, 0.00019292, 
    0.00018692, 0.00018111, 0.00017532, 0.00016964, 0.00016428, 0.0001592, 
    0.00015442, 0.00014973, 0.00014508, 0.0001405, 0.00013602, 0.00013179, 
    0.00012765, 0.00012352, 0.00011954, 0.00011551, 0.00011145, 0.00010744, 
    0.00010347, 9.963e-05, 9.59e-05, 9.246e-05, 8.933e-05, 8.623e-05, 
    8.324e-05, 8.001e-05, 7.678e-05, 7.361e-05, 7.075e-05, 6.834e-05, 
    6.628e-05, 6.443e-05, 6.246e-05, 6.042e-05, 5.822e-05, 5.602e-05, 
    5.406e-05, 5.229e-05, 5.08e-05, 4.93e-05, 4.786e-05, 4.645e-05, 
    4.508e-05, 4.371e-05, 4.229e-05, 4.091e-05, 3.951e-05, 3.813e-05, 
    3.692e-05, 3.572e-05, 3.451e-05, 3.331e-05, 3.234e-05, 3.157e-05, 
    3.072e-05, 2.964e-05, 2.852e-05, 2.755e-05, 2.668e-05, 2.59e-05, 
    2.522e-05, 2.489e-05, 2.473e-05, 2.434e-05, 2.298e-05, 2.049e-05, 
    1.825e-05, 1.753e-05, 1.866e-05, 2.031e-05, 2.045e-05, 1.967e-05, 
    1.88e-05, 1.841e-05, 1.857e-05, 1.849e-05, 1.771e-05, 1.628e-05, 
    1.489e-05, 1.406e-05, 1.385e-05, 1.376e-05, 1.366e-05, 1.344e-05, 
    1.326e-05, 1.314e-05, 1.294e-05, 1.258e-05, 1.238e-05, 1.181e-05, 
    1.116e-05, 1.073e-05, 1.034e-05, 9.83e-06, 9.25e-06, 8.85e-06, 8.54e-06, 
    8.24e-06, 7.83e-06, 7.64e-06, 7.79e-06, 8.15e-06, 8.77e-06, 9.5e-06, 
    9.54e-06, 8.91e-06, 8.2e-06, 7.69e-06, 7.52e-06, 7.48e-06, 7.33e-06, 
    6.69e-06, 5.91e-06, 5.2e-06, 4.77e-06, 4.52e-06, 4.3e-06, 4.13e-06, 
    4.53e-06, 5.51e-06, 6.18e-06, 6.26e-06, 5.36e-06, 3.61e-06, 2.05e-06, 
    1.54e-06, 2.47e-06, 3.42e-06, 3.88e-06, 3.98e-06, 3.81e-06, 4.15e-06, 
    4.67e-06, 4.79e-06, 4.54e-06, 3.95e-06, 3.36e-06, 3.08e-06, 2.99e-06, 
    3.05e-06, 2.76e-06, 2.74e-06, 3.1e-06, 3.84e-06, 4.46e-06, 4.38e-06, 
    3.96e-06, 3.59e-06, 3.26e-06, 2.91e-06, 2.46e-06, 2.23e-06, 2.35e-06, 
    2.55e-06, 2.85e-06, 3.82e-06, 4.01e-06, 3.37e-06, 2.5e-06, 2.05e-06, 
    1.91e-06, 1.82e-06, 1.75e-06, 1.68e-06, 1.8e-06, 2.17e-06, 2.48e-06, 
    2.7e-06, 2.85e-06, 2.96e-06, 2.75e-06, 2.32e-06, 1.85e-06, 1.55e-06, 
    1.44e-06, 1.26e-06, 8.9e-07, 7.3e-07, 7.9e-07, 9.4e-07, 8.2e-07, 7.1e-07, 
    6.7e-07, 6.9e-07, 8.7e-07, 1.22e-06, 1.76e-06, 2.05e-06, 1.82e-06, 
    1.2e-06, 6.8e-07, 4.8e-07, 3.6e-07, 1.5e-07, 2e-07, 2.1e-07, 1.3e-07, 
    -2.4e-07, -6.2e-07, 4e-08, 1.16e-06, 2.07e-06, 2.11e-06 ;

 bangle_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 alt_refrac =
  18263, 18571, 18879, 19186, 19494, 19800, 20106, 20411, 20716, 21022, 
    21327, 21631, 21936, 22240, 22544, 22848, 23152, 23455, 23759, 24062, 
    24365, 24669, 24972, 25274, 25576, 25879, 26181, 26483, 26785, 27086, 
    27388, 27690, 27991, 28293, 28594, 28896, 29197, 29498, 29799, 30100, 
    30401, 30702, 31003, 31304, 31605, 31906, 32207, 32507, 32808, 33108, 
    33409, 33710, 34010, 34310, 34611, 34911, 35212, 35512, 35812, 36113, 
    36413, 36713, 37014, 37314, 37614, 37914, 38214, 38515, 38815, 39115, 
    39415, 39715, 40015, 40315, 40615, 40915, 41215, 41515, 41815, 42115, 
    42415, 42715, 43015, 43315, 43615, 43915, 44215, 44515, 44815, 45115, 
    45415, 45715, 46014, 46314, 46614, 46914, 47214, 47514, 47814, 48114, 
    48414, 48714, 49013, 49313, 49613, 49913, 50213, 50513, 50813, 51112, 
    51412, 51712, 52012, 52312, 52612, 52911, 53211, 53511, 53811, 54111, 
    54411, 54711, 55010, 55310, 55610, 55910, 56210, 56509, 56809, 57109, 
    57409, 57709, 58009, 58308, 58608, 58908, 59208, 59508, 59808, 60107, 
    60407, 60707, 61007, 61307, 61606, 61906, 62206, 62506, 62806, 63105, 
    63405, 63705, 64005, 64305, 64605, 64904, 65204, 65504, 65804, 66104, 
    66403, 66703, 67003, 67303, 67603, 67902, 68202, 68502, 68802, 69102, 
    69401, 69701, 70001, 70301, 70601, 70900, 71200, 71500, 71800, 72100, 
    72399, 72699, 72999, 73299, 73599, 73899, 74198, 74498, 74798, 75098, 
    75398, 75697, 75997, 76297, 76597, 76897, 77196, 77496, 77796, 78096, 
    78396, 78695, 78995, 79295, 79595, 79895, 80194, 80494, 80794, 81094, 
    81394, 81693, 81993, 82293, 82593, 82893, 83192, 83492, 83792, 84092, 
    84392, 84691, 84991, 85291, 85591, 85891, 86190, 86490, 86790, 87090, 
    87390, 87689, 87989, 88289, 88589, 88889, 89188, 89488, 89788, 90088, 
    90388, 90687, 90987, 91287, 91587, 91887, 92186, 92486, 92786, 93086, 
    93386, 93685, 93985, 94285, 94585, 94885, 95184, 95484, 95784, 96084, 
    96383, 96683, 96983, 97283, 97583, 97882, 98182, 98482, 98782, 99082, 
    99381, 99681, 99981 ;

 geop_refrac =
  18219, 18525, 18832, 19137, 19443, 19748, 20052, 20355, 20658, 20962, 
    21266, 21568, 21871, 22173, 22475, 22777, 23079, 23380, 23682, 23982, 
    24283, 24585, 24886, 25186, 25485, 25786, 26086, 26385, 26685, 26984, 
    27283, 27583, 27881, 28181, 28479, 28779, 29077, 29375, 29674, 29972, 
    30270, 30569, 30867, 31165, 31463, 31761, 32060, 32357, 32655, 32952, 
    33250, 33548, 33845, 34142, 34440, 34736, 35034, 35331, 35628, 35926, 
    36222, 36519, 36817, 37114, 37410, 37707, 38003, 38301, 38597, 38894, 
    39190, 39487, 39783, 40080, 40376, 40672, 40969, 41265, 41561, 41857, 
    42154, 42450, 42746, 43042, 43338, 43634, 43930, 44226, 44522, 44818, 
    45114, 45410, 45705, 46000, 46296, 46592, 46888, 47183, 47479, 47775, 
    48070, 48366, 48661, 48956, 49252, 49547, 49843, 50138, 50434, 50728, 
    51023, 51319, 51614, 51909, 52204, 52499, 52794, 53089, 53384, 53679, 
    53974, 54269, 54564, 54859, 55153, 55448, 55743, 56037, 56332, 56627, 
    56922, 57217, 57511, 57805, 58100, 58394, 58689, 58984, 59278, 59572, 
    59866, 60161, 60455, 60750, 61043, 61338, 61632, 61926, 62221, 62514, 
    62808, 63102, 63397, 63691, 63985, 64278, 64572, 64866, 65160, 65454, 
    65747, 66041, 66335, 66629, 66923, 67216, 67510, 67803, 68097, 68391, 
    68684, 68977, 69271, 69565, 69858, 70151, 70444, 70738, 71031, 71325, 
    71617, 71911, 72204, 72497, 72791, 73084, 73376, 73670, 73963, 74256, 
    74549, 74841, 75134, 75427, 75721, 76014, 76306, 76599, 76891, 77184, 
    77477, 77769, 78062, 78355, 78648, 78940, 79232, 79525, 79817, 80110, 
    80403, 80694, 80987, 81279, 81572, 81864, 82156, 82448, 82741, 83033, 
    83325, 83617, 83909, 84201, 84494, 84786, 85077, 85369, 85661, 85953, 
    86245, 86536, 86828, 87120, 87412, 87704, 87995, 88287, 88579, 88871, 
    89163, 89453, 89745, 90037, 90329, 90620, 90911, 91203, 91494, 91786, 
    92077, 92368, 92659, 92951, 93242, 93534, 93824, 94115, 94407, 94698, 
    94988, 95279, 95571, 95862, 96153, 96443, 96734, 97025, 97316, 97607, 
    97897, 98188, 98479 ;

 refrac =
  27.079, 25.788, 24.527, 23.283, 22.119, 21.11, 20.186, 19.292, 18.419, 
    17.575, 16.765, 16.007, 15.273, 14.544, 13.842, 13.196, 12.608, 12.051, 
    11.495, 10.927, 10.364, 9.833, 9.351, 8.917, 8.516, 8.138, 7.779, 7.438, 
    7.113, 6.801, 6.5, 6.21, 5.93, 5.66, 5.399, 5.152, 4.921, 4.706, 4.501, 
    4.303, 4.113, 3.931, 3.757, 3.589, 3.425, 3.268, 3.118, 2.977, 2.845, 
    2.723, 2.609, 2.498, 2.39, 2.286, 2.188, 2.095, 2.006, 1.919, 1.836, 
    1.755, 1.678, 1.604, 1.533, 1.464, 1.398, 1.335, 1.275, 1.218, 1.164, 
    1.113, 1.064, 1.017, 0.974, 0.935, 0.899, 0.864, 0.828, 0.793, 0.76, 
    0.729, 0.7, 0.673, 0.647, 0.622, 0.598, 0.574, 0.551, 0.53, 0.51, 0.491, 
    0.472, 0.453, 0.436, 0.421, 0.405, 0.388, 0.374, 0.363, 0.352, 0.338, 
    0.321, 0.307, 0.298, 0.289, 0.28, 0.271, 0.262, 0.253, 0.243, 0.233, 
    0.224, 0.215, 0.207, 0.199, 0.193, 0.187, 0.18, 0.173, 0.167, 0.161, 
    0.155, 0.149, 0.143, 0.138, 0.133, 0.129, 0.124, 0.12, 0.116, 0.113, 
    0.109, 0.105, 0.1, 0.097, 0.093, 0.09, 0.086, 0.083, 0.08, 0.077, 0.074, 
    0.072, 0.069, 0.066, 0.064, 0.061, 0.059, 0.056, 0.054, 0.053, 0.051, 
    0.049, 0.047, 0.045, 0.043, 0.042, 0.04, 0.038, 0.037, 0.035, 0.034, 
    0.033, 0.031, 0.03, 0.029, 0.028, 0.026, 0.025, 0.024, 0.023, 0.022, 
    0.021, 0.021, 0.02, 0.019, 0.018, 0.017, 0.017, 0.016, 0.015, 0.015, 
    0.014, 0.013, 0.013, 0.012, 0.012, 0.011, 0.011, 0.01, 0.01, 0.009, 
    0.009, 0.009, 0.008, 0.008, 0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 
    0.006, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 refrac_sigma =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 refrac_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 dry_temp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 dry_temp_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 dry_temp_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;
}
