netcdf ropp_test_2v {
dimensions:
	dim_unlim = UNLIMITED ; // (1 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1a = 100 ;
	dim_lev1b = 100 ;
	dim_lev2a = 100 ;
	dim_lev2b = 100 ;
	dim_lev2d = 100 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 360. ;
	char bg_source(dim_unlim, dim_char20) ;
		bg_source:long_name = "Background data source" ;
	int bg_year(dim_unlim) ;
		bg_year:long_name = "VT year" ;
		bg_year:units = "years" ;
		bg_year:valid_range = 1995, 2099 ;
	int bg_month(dim_unlim) ;
		bg_month:long_name = "VT month" ;
		bg_month:units = "months" ;
		bg_month:valid_range = 1, 12 ;
	int bg_day(dim_unlim) ;
		bg_day:long_name = "VT day" ;
		bg_day:units = "days" ;
		bg_day:valid_range = 1, 31 ;
	int bg_hour(dim_unlim) ;
		bg_hour:long_name = "VT hour" ;
		bg_hour:units = "hours" ;
		bg_hour:valid_range = 0, 23 ;
	int bg_minute(dim_unlim) ;
		bg_minute:long_name = "VT minute" ;
		bg_minute:units = "minutes" ;
		bg_minute:valid_range = 0, 59 ;
	float bg_fcperiod(dim_unlim) ;
		bg_fcperiod:long_name = "Forecast period" ;
		bg_fcperiod:units = "hours" ;
		bg_fcperiod:valid_range = 0., 24. ;
	double dtime(dim_unlim, dim_lev1a) ;
		dtime:long_name = "Time since start of occultation" ;
		dtime:units = "seconds" ;
		dtime:valid_range = -1., 240. ;
	float snr_L1ca(dim_unlim, dim_lev1a) ;
		snr_L1ca:long_name = "Signal-to-noise ratio (L1, C/A code)" ;
		snr_L1ca:units = "volt / volt" ;
		snr_L1ca:valid_range = 0., 50000. ;
	float snr_L1p(dim_unlim, dim_lev1a) ;
		snr_L1p:long_name = "Signal-to-noise ratio (L1, P code)" ;
		snr_L1p:units = "volt / volt" ;
		snr_L1p:valid_range = 0., 50000. ;
	float snr_L2p(dim_unlim, dim_lev1a) ;
		snr_L2p:long_name = "Signal-to-noise ratio (L2, P code)" ;
		snr_L2p:units = "volt / volt" ;
		snr_L2p:valid_range = 0., 50000. ;
	double phase_L1(dim_unlim, dim_lev1a) ;
		phase_L1:long_name = "Excess phase (L1)" ;
		phase_L1:units = "metres" ;
		phase_L1:valid_range = -1.e+06, 1.e+06 ;
	double phase_L2(dim_unlim, dim_lev1a) ;
		phase_L2:long_name = "Excess phase (L2)" ;
		phase_L2:units = "metres" ;
		phase_L2:valid_range = -1.e+06, 1.e+06 ;
	double r_gns(dim_unlim, xyz, dim_lev1a) ;
		r_gns:long_name = "GNSS transmitter position" ;
		r_gns:units = "metres" ;
		r_gns:valid_range = -4.3e+07, 4.3e+07 ;
		r_gns:reference_frame = "ECF" ;
	double v_gns(dim_unlim, xyz, dim_lev1a) ;
		v_gns:long_name = "GNSS transmitter velocity" ;
		v_gns:units = "metres / seconds" ;
		v_gns:valid_range = -10000., 10000. ;
		v_gns:reference_frame = "ECI" ;
	double r_leo(dim_unlim, xyz, dim_lev1a) ;
		r_leo:long_name = "LEO transmitter position" ;
		r_leo:units = "metres" ;
		r_leo:valid_range = -1.e+07, 1.e+07 ;
		r_leo:reference_frame = "ECF" ;
	double v_leo(dim_unlim, xyz, dim_lev1a) ;
		v_leo:long_name = "LEO transmitter velocity" ;
		v_leo:units = "metres / seconds" ;
		v_leo:valid_range = -10000., 10000. ;
		v_leo:reference_frame = "ECI" ;
	float phase_qual(dim_unlim, dim_lev1a) ;
		phase_qual:long_name = "Quality value for phase (and SNR)" ;
		phase_qual:units = "percent" ;
		phase_qual:valid_range = 0., 100. ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 360. ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float alt_refrac(dim_unlim, dim_lev2a) ;
		alt_refrac:long_name = "Geometric height above geoid for refractivity" ;
		alt_refrac:units = "metres" ;
		alt_refrac:valid_range = -1000., 1.e+05 ;
	float geop_refrac(dim_unlim, dim_lev2a) ;
		geop_refrac:long_name = "Geopotential height above geoid for refractivity" ;
		geop_refrac:units = "geopotential metres" ;
		geop_refrac:valid_range = -1000., 1.e+05 ;
	double refrac(dim_unlim, dim_lev2a) ;
		refrac:long_name = "Refractivity" ;
		refrac:units = "N-units" ;
		refrac:valid_range = 0., 500. ;
	double refrac_sigma(dim_unlim, dim_lev2a) ;
		refrac_sigma:long_name = "Estimated error (1-sigma) for refractivity" ;
		refrac_sigma:units = "N-units" ;
		refrac_sigma:valid_range = 0., 50. ;
	float refrac_qual(dim_unlim, dim_lev2a) ;
		refrac_qual:long_name = "Quality value for refractivity" ;
		refrac_qual:units = "percent" ;
		refrac_qual:valid_range = 0., 100. ;
	double dry_temp(dim_unlim, dim_lev2a) ;
		dry_temp:long_name = "Dry temperature" ;
		dry_temp:units = "kelvin" ;
		dry_temp:valid_range = 150., 350. ;
	double dry_temp_sigma(dim_unlim, dim_lev2a) ;
		dry_temp_sigma:long_name = "Estimated error (1-sigma) for dry temperature" ;
		dry_temp_sigma:units = "kelvin" ;
		dry_temp_sigma:valid_range = 0., 50. ;
	float dry_temp_qual(dim_unlim, dim_lev2a) ;
		dry_temp_qual:long_name = "Quality value for dry temperature" ;
		dry_temp_qual:units = "percent" ;
		dry_temp_qual:valid_range = 0., 100. ;
	float geop(dim_unlim, dim_lev2b) ;
		geop:long_name = "Geopotential height above geoid for P,T,H" ;
		geop:units = "geopotential metres" ;
		geop:valid_range = -1000., 1.e+05 ;
	float geop_sigma(dim_unlim, dim_lev2b) ;
		geop_sigma:long_name = "Estimated error (1-sigma) for geopotential height" ;
		geop_sigma:units = "geopotential metres" ;
		geop_sigma:valid_range = 0., 500. ;
	double press(dim_unlim, dim_lev2b) ;
		press:long_name = "Pressure" ;
		press:units = "hPa" ;
		press:valid_range = 0.0001, 1100. ;
	float press_sigma(dim_unlim, dim_lev2b) ;
		press_sigma:long_name = "Estimated error (1-sigma) for pressure" ;
		press_sigma:units = "hPa" ;
		press_sigma:valid_range = 0., 5. ;
	double temp(dim_unlim, dim_lev2b) ;
		temp:long_name = "Temperature" ;
		temp:units = "kelvin" ;
		temp:valid_range = 150., 350. ;
	float temp_sigma(dim_unlim, dim_lev2b) ;
		temp_sigma:long_name = "Estimated error (1-sigma) for temperature" ;
		temp_sigma:units = "kelvin" ;
		temp_sigma:valid_range = 0., 5. ;
	double shum(dim_unlim, dim_lev2b) ;
		shum:long_name = "Specific humidity" ;
		shum:units = "gram / kilogram" ;
		shum:valid_range = 0., 50. ;
	float shum_sigma(dim_unlim, dim_lev2b) ;
		shum_sigma:long_name = "Estimated  error (1-sigma) in specific humidity" ;
		shum_sigma:units = "gram / kilogram" ;
		shum_sigma:valid_range = 0., 5. ;
	float meteo_qual(dim_unlim, dim_lev2b) ;
		meteo_qual:long_name = "Quality value for meteorological data" ;
		meteo_qual:units = "percent" ;
		meteo_qual:valid_range = 0., 100. ;
	float geop_sfc(dim_unlim) ;
		geop_sfc:long_name = "Surface geopotential height" ;
		geop_sfc:units = "geopotential metres" ;
		geop_sfc:valid_range = -1000., 10000. ;
	float press_sfc(dim_unlim) ;
		press_sfc:long_name = "Surface pressure" ;
		press_sfc:units = "hPa" ;
		press_sfc:valid_range = 250., 1100. ;
	float press_sfc_sigma(dim_unlim) ;
		press_sfc_sigma:long_name = "Estimated error (1-sigma) for surface pressure" ;
		press_sfc_sigma:units = "hPa" ;
		press_sfc_sigma:valid_range = 0., 5. ;
	float press_sfc_qual(dim_unlim) ;
		press_sfc_qual:long_name = "Surface pressure quality value" ;
		press_sfc_qual:units = "percent" ;
		press_sfc_qual:valid_range = 0., 100. ;
	double tph_bangle(dim_unlim) ;
		tph_bangle:long_name = "Bending angle-based TPH" ;
		tph_bangle:units = "metres" ;
		tph_bangle:valid_range = 6.2e+06, 6.6e+06 ;
	double tpa_bangle(dim_unlim) ;
		tpa_bangle:long_name = "Bending angle-based TPA" ;
		tpa_bangle:units = "radians" ;
		tpa_bangle:valid_range = -0.001, 0.1 ;
	int tph_bangle_flag(dim_unlim) ;
		tph_bangle_flag:long_name = "Bending angle-based TPH QC flag" ;
		tph_bangle_flag:units = "1" ;
		tph_bangle_flag:valid_range = 0, 255 ;
	float tph_refrac(dim_unlim) ;
		tph_refrac:long_name = "Refractivity-based TPH" ;
		tph_refrac:units = "metres" ;
		tph_refrac:valid_range = -1000., 1.e+05 ;
	double tpn_refrac(dim_unlim) ;
		tpn_refrac:long_name = "Refractivity-based TPN" ;
		tpn_refrac:units = "N-units" ;
		tpn_refrac:valid_range = 0., 500. ;
	int tph_refrac_flag(dim_unlim) ;
		tph_refrac_flag:long_name = "Refractivity-based TPH QC flag" ;
		tph_refrac_flag:units = "1" ;
		tph_refrac_flag:valid_range = 0, 255 ;
	float tph_tdry_lrt(dim_unlim) ;
		tph_tdry_lrt:long_name = "Dry temperature-based TPH (lapse rate)" ;
		tph_tdry_lrt:units = "metres" ;
		tph_tdry_lrt:valid_range = -1000., 1.e+05 ;
	float tpt_tdry_lrt(dim_unlim) ;
		tpt_tdry_lrt:long_name = "Dry temperature-based TPT (lapse rate)" ;
		tpt_tdry_lrt:units = "kelvin" ;
		tpt_tdry_lrt:valid_range = 150., 350. ;
	int tph_tdry_lrt_flag(dim_unlim) ;
		tph_tdry_lrt_flag:long_name = "Dry temperature-based TPH QC flag (lapse rate)" ;
		tph_tdry_lrt_flag:units = "1" ;
		tph_tdry_lrt_flag:valid_range = 0, 255 ;
	float tph_tdry_cpt(dim_unlim) ;
		tph_tdry_cpt:long_name = "Dry temperature-based TPH (cold point)" ;
		tph_tdry_cpt:units = "metres" ;
		tph_tdry_cpt:valid_range = -1000., 1.e+05 ;
	float tpt_tdry_cpt(dim_unlim) ;
		tpt_tdry_cpt:long_name = "Dry temperature-based TPT (cold point)" ;
		tpt_tdry_cpt:units = "kelvin" ;
		tpt_tdry_cpt:valid_range = 150., 350. ;
	int tph_tdry_cpt_flag(dim_unlim) ;
		tph_tdry_cpt_flag:long_name = "Dry temperature-based TPH QC flag (cold point)" ;
		tph_tdry_cpt_flag:units = "1" ;
		tph_tdry_cpt_flag:valid_range = 0, 255 ;
	float prh_tdry_cpt(dim_unlim) ;
		prh_tdry_cpt:long_name = "Dry temperature-based PRH (cold point)" ;
		prh_tdry_cpt:units = "metres" ;
	float prt_tdry_cpt(dim_unlim) ;
		prt_tdry_cpt:long_name = "Dry temperature-based PRT (cold point)" ;
		prt_tdry_cpt:units = "kelvin" ;
	int prh_tdry_cpt_flag(dim_unlim) ;
		prh_tdry_cpt_flag:long_name = "Dry temperature-based PRH QC flag (cold point)" ;
		prh_tdry_cpt_flag:units = "1" ;
	float tph_temp_lrt(dim_unlim) ;
		tph_temp_lrt:long_name = "Temperature-based TPH (lapse rate)" ;
		tph_temp_lrt:units = "geopotential metres" ;
		tph_temp_lrt:valid_range = -1000., 1.e+05 ;
	float tpt_temp_lrt(dim_unlim) ;
		tpt_temp_lrt:long_name = "Temperature-based TPT (lapse rate)" ;
		tpt_temp_lrt:units = "kelvin" ;
		tpt_temp_lrt:valid_range = 150., 350. ;
	int tph_temp_lrt_flag(dim_unlim) ;
		tph_temp_lrt_flag:long_name = "Temperature-based TPH QC flag (lapse rate)" ;
		tph_temp_lrt_flag:units = "1" ;
		tph_temp_lrt_flag:valid_range = 0, 255 ;
	float tph_temp_cpt(dim_unlim) ;
		tph_temp_cpt:long_name = "Temperature-based TPH (cold point)" ;
		tph_temp_cpt:units = "geopotential metres" ;
		tph_temp_cpt:valid_range = -1000., 1.e+05 ;
	float tpt_temp_cpt(dim_unlim) ;
		tpt_temp_cpt:long_name = "Temperature-based TPT (cold point)" ;
		tpt_temp_cpt:units = "kelvin" ;
		tpt_temp_cpt:valid_range = 150., 350. ;
	int tph_temp_cpt_flag(dim_unlim) ;
		tph_temp_cpt_flag:long_name = "Temperature-based TPH QC flag (cold point)" ;
		tph_temp_cpt_flag:units = "1" ;
		tph_temp_cpt_flag:valid_range = 0, 255 ;
	float prh_temp_cpt(dim_unlim) ;
		prh_temp_cpt:long_name = "Temperature-based PRH (cold point)" ;
		prh_temp_cpt:units = "metres" ;
	float prt_temp_cpt(dim_unlim) ;
		prt_temp_cpt:long_name = "Temperature-based PRT (cold point)" ;
		prt_temp_cpt:units = "kelvin" ;
	int prh_temp_cpt_flag(dim_unlim) ;
		prh_temp_cpt_flag:long_name = "Temperature-based PRH QC flag (cold point)" ;
		prh_temp_cpt_flag:units = "1" ;
	char level_type(dim_unlim, dim_char64) ;
		level_type:long_name = "Vertical level type" ;
	float level_coeff_a(dim_unlim, dim_lev2d) ;
		level_coeff_a:long_name = "Hybrid / Eta level coefficient (a or eta)" ;
		level_coeff_a:units = "hPa" ;
		level_coeff_a:valid_range = 0., 2000. ;
	float level_coeff_b(dim_unlim, dim_lev2d) ;
		level_coeff_b:long_name = "Hybrid / Eta level coefficient (b or tau)" ;
		level_coeff_b:units = "1" ;
		level_coeff_b:valid_range = 0., 2. ;

// global attributes:
		:title = "Atmospheric background data for ROPP Radio Occultation data" ;
		:institution = "HIRLAM" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "NESDIS" ;
		:processing_date = "2014-11-26 10:20:25.893" ;
		:pod_method = "POD_5" ;
		:phase_method = "PHASE_2" ;
		:bangle_method = "BANGLE_4" ;
		:refrac_method = "REFRAC_6" ;
		:meteo_method = "T-DRY" ;
		:thin_method = "ASGLIN" ;
		:software_version = "V35.348" ;
		:_FillValue = -9.9999e+07 ;
data:

 occ_id =
  "BG_20141028001753_CHMP_R016_NESD" ;

 gns_id =
  "R016" ;

 leo_id =
  "CHMP" ;

 stn_id =
  "KIRU" ;

 start_time = 4.6777e+08 ;

 year = 2014 ;

 month = 10 ;

 day = 28 ;

 hour = 0 ;

 minute = 17 ;

 second = 53 ;

 msec = 46 ;

 pcd = 19089 ;

 overall_qual = 92.098 ;

 time = 4.6777e+08 ;

 time_offset = 174.96 ;

 lat = 34.929 ;

 lon = 45.02 ;

 undulation = -68.868 ;

 roc = 6.2568e+06 ;

 r_coc =
  19970, 5987, -34689 ;

 azimuth = 23.973 ;

 bg_source =
  "HIRLAM" ;

 bg_year = 2014 ;

 bg_month = 10 ;

 bg_day = 28 ;

 bg_hour = 18 ;

 bg_minute = 0 ;

 bg_fcperiod = 3 ;

 dtime =
  52.036, 26.654, 18.151, -0.8665, 31.944, 108.9, 191.35, 130.33, 192.91, 
    24.485, 35.694, 193.25, 123.99, 39.544, 200.76, 87.602, 19.131, 155.73, 
    145.05, 14.854, 194.04, 183.8, 144.48, 50.009, 128.39, 128.21, 191.79, 
    219.64, 68.105, 29.567, 223.32, 70.745, 55.11, 152.81, 25.315, 209.45, 
    25.885, 132.08, 158.13, 64.788, 119.59, 177.02, 23.201, 151.58, -0.77278, 
    19.111, 60.92, 186.16, 11.366, 2.4487, 16.604, 141.71, 232.53, 83.053, 
    66.859, 35.575, 115.97, 133.37, 130.18, 111.56, 154.85, 67.25, 227.27, 
    49.305, 122.08, 78.368, 138.68, 43.789, 214.89, 99.659, 1.6124, 177.72, 
    116.68, 163.79, 78.74, 132.73, 73.44, 41.129, 97.082, 63.528, 107.97, 
    206.17, 225.85, 81.993, 69.436, 95.408, 173.72, 233.81, 139.03, 119.79, 
    204, 191.51, 218, 118.2, 90.55, 44.226, 46.081, 46.929, 27.636, 194.6 ;

 snr_L1ca =
  35170, 28978, 28840, 35864, 32337, 42820, 47756, 41109, 41284, 26596, 
    29433, 36179, 15322, 38687, 26881, 22728, 44703, 1618.5, 2784.2, 66.777, 
    676.61, 21347, 12140, 11295, 2161.3, 20986, 39616, 8877.3, 21330, 25036, 
    17893, 36522, 2765.9, 10301, 10459, 20986, 779.68, 46876, 32476, 44470, 
    26755, 41704, 13593, 18499, 47224, 13437, 30664, 20486, 17649, 32060, 
    32857, 5927.4, 11169, 20785, 15404, 26187, 40624, 21436, 22604, 63.887, 
    3881.6, 7630.3, 32278, 41805, 16733, 4995.8, 30418, 33475, 9497.4, 47522, 
    20450, 42105, 14186, 35982, 28989, 15248, 5733.7, 32183, 34705, 12537, 
    37671, 36336, 27094, 11741, 23173, 45711, 47470, 41605, 34550, 30897, 
    27522, 30253, 44671, 45060, 46111, 45959, 4438.3, 21542, 45.025, 23878 ;

 snr_L1p =
  47601, 47874, 19657, 19338, 11231, 42239, 36635, 7011.8, 14081, 16742, 
    46304, 33994, 42877, 7952.7, 32746, 905.22, 26501, 20321, 31778, 13448, 
    18909, 11885, 21497, 29121, 23309, 21097, 46989, 23801, 13322, 39842, 
    25469, 32215, 48102, 37457, 38636, 29138, 37959, 37736, 20467, 14467, 
    43612, 6669.8, 3150.3, 5978.8, 29065, 18480, 47862, 45564, 22205, 8131.7, 
    46850, 22889, 6374, 24606, 25539, 555.52, 17617, 18921, 28374, 37120, 
    29869, 48991, 13506, 4078.9, 46147, 5861.8, 23613, 33510, 33097, 19707, 
    37154, 19546, 38282, 4900.6, 22355, 47946, 36773, 11787, 2686.7, 8537.8, 
    23725, 3984.7, 39877, 27152, 30240, 5595.3, 7547.5, 18371, 35897, 7191.5, 
    32828, 17266, 31478, 4266.5, 20856, 35426, 8301.4, 3454.3, 47542, 11982 ;

 snr_L2p =
  45210, 42346, 27607, 17418, 8474.8, 27838, 13603, 18896, 6616.9, 14797, 
    20305, 447.12, 44334, 45463, 16852, 45983, 20027, 14624, 35085, 31654, 
    18832, 48640, 40021, 45742, 24095, 25428, 7148.9, 11950, 23494, 20401, 
    19851, 13353, 199.24, 20296, 37093, 11175, 48696, 23863, 45830, 35721, 
    7116.6, 32055, 8772.1, 30595, 30983, 32147, 46809, 5665.7, 41031, 20763, 
    29659, 15765, 37633, 34717, 17559, 12060, 23532, 5164.5, 5408.7, 24755, 
    43206, 20220, 31861, 46027, 37989, 47347, 9892.4, 5651.9, 17631, 46917, 
    23582, 21414, 13126, 39217, 8399.2, 11988, 47660, 11523, 6952.3, 8876.8, 
    12432, 35496, 35447, 43637, 8578.3, 28362, 44324, 41727, 9169.3, 41381, 
    34966, 6969.3, 16275, 42872, 36550, 20296, 760.03, 2365, 27554, 47468 ;

 phase_L1 =
  -6.4712e+05, -2.7874e+05, 2.2615e+05, 8.4768e+05, -3.3919e+05, -8.6841e+05, 
    9.405e+05, 1.8752e+05, -9.1961e+05, 743.75, 67656, 6.2883e+05, 
    9.3043e+05, 3.8752e+05, -3.5157e+05, 3.2985e+05, -7.9152e+05, -59073, 
    6.9521e+05, -2.7908e+05, -3.1094e+05, 1.3504e+05, -2.7983e+05, 
    -3.8292e+05, -8.8075e+05, -8.2922e+05, 6.4859e+05, 8.9389e+05, 
    -8.9304e+05, 6.323e+05, -4.6905e+05, 8.6999e+05, 3.5782e+05, 1.9746e+05, 
    1.3234e+05, -5.5411e+05, 3.6465e+05, 8.3342e+05, 8.6008e+05, 15587, 
    -1.4622e+05, 58903, 5.3821e+05, -67831, -8.786e+05, 2.1934e+05, 
    -8.4413e+05, 6.074e+05, -6.4292e+05, -73537, -3.9384e+05, 4.4416e+05, 
    -7.2544e+05, -9.9846e+05, 8.5352e+05, -7.1541e+05, -4.5674e+05, 
    -9.8297e+05, -96934, -68528, -2.7687e+05, -7.4928e+05, 1.3566e+05, 
    6.836e+05, 1.4561e+05, -4.4103e+05, -27596, -2.7208e+05, 9.2955e+05, 
    -4.279e+05, 6.1148e+05, -6.8207e+05, -2.2986e+05, -7.8134e+05, 
    6.7542e+05, 6.6735e+05, -2.7268e+05, 4.7049e+05, -8.4953e+05, 
    -5.5621e+05, 4.809e+05, -4.2809e+05, -20825, 7.5193e+05, -9.461e+05, 
    6.6933e+05, 9.1372e+05, -4.6737e+05, 1.6521e+05, -9.5991e+05, 
    -8.9628e+05, -5.2279e+05, -87170, 67762, 7.3044e+05, 5.2504e+05, 
    7.6445e+05, -9.5879e+05, -70188, 3.4668e+05 ;

 phase_L2 =
  1.5788e+05, -47156, -1.9819e+05, -2.4657e+05, -5.3945e+05, -5.0691e+05, 
    1.3505e+05, -11039, -8.7036e+05, 45690, -2.9291e+05, 5.688e+05, 
    -2.9888e+05, 6.3689e+05, 5.866e+05, 9.5598e+05, -8.1446e+05, -4.5778e+05, 
    -8.6218e+05, 1.3087e+05, -4.3127e+05, -84233, -8.4566e+05, 3.6158e+05, 
    3.1479e+05, 2.7788e+05, -6.4798e+05, -5.185e+05, -8.2493e+05, 
    -6.6817e+05, 5.6026e+05, 1.3511e+05, -7.8321e+05, -2.0617e+05, 
    7.1522e+05, 57734, 4.6309e+05, 3.9559e+05, -5.3606e+05, 6.8923e+05, 
    -4.4534e+05, 3.2943e+05, -5.7455e+05, 7.5608e+05, 5.2913e+05, 
    -6.9652e+05, -5.2215e+05, 8.9935e+05, -5.6483e+05, 8.8474e+05, 
    2.6035e+05, -1.8141e+05, -1.7222e+05, -6.7892e+05, -7.288e+05, 
    5.4666e+05, -7.6021e+05, 6.5225e+05, 4.8241e+05, 5.3695e+05, 7.3177e+05, 
    7.156e+05, -4.0234e+05, -7.538e+05, -5.7703e+05, -6.4211e+05, -7.633e+05, 
    5.9872e+05, -8.5244e+05, 3.7598e+05, -4.4042e+05, 6.517e+05, -1.0682e+05, 
    8.3943e+05, -1.8584e+05, -7.222e+05, 6.7987e+05, 8.6073e+05, -4.4655e+05, 
    1.5851e+05, 7.063e+05, 36496, 9.5288e+05, -7.0322e+05, -4.3545e+05, 
    7.8579e+05, -7.3754e+05, 8.2093e+05, 1.5179e+05, -3.2643e+05, 
    -5.2297e+05, 19757, 2.4222e+05, -8.9917e+05, -7.4456e+05, -9.4762e+05, 
    1.1773e+05, -9.5686e+05, 36246, 3.6398e+05 ;

 r_gns =
  4.1918e+06, -2.2774e+07, -4.9857e+06, 4.9093e+06, -3.4331e+06, -8.9421e+06, 
    -1.9681e+05, -1.0605e+07, 4.0878e+06, 2.1651e+07, 3.1488e+06, 2.4826e+07, 
    5.3112e+06, -4.7562e+06, 1.3494e+05, -1.1739e+07, 1.0584e+07, 1.4743e+07, 
    6.7242e+06, 1.7731e+07, 2.0272e+07, -8.3863e+06, -9.5053e+05, 
    -9.9204e+05, 4.9099e+06, 7.2277e+05, 9.4284e+06, 2.8521e+07, 2.387e+05, 
    -9.0096e+06, -4.4334e+05, -1.6376e+06, -1.2409e+06, 6.4848e+06, 
    -7.9067e+05, 3.9839e+06, 1.1126e+07, 4.8844e+06, -1.8836e+06, 
    -1.4154e+07, 2.3087e+07, 3.0782e+06, -1.3759e+07, 5.2362e+06, 9.8255e+05, 
    1.132e+07, 2.72e+07, -9.2202e+06, 1.0689e+07, 9.1676e+06, -3.1242e+06, 
    -1.05e+07, 3.0861e+06, -1.1234e+06, -1.0508e+07, 2.339e+06, 4.8787e+06, 
    -8.8438e+06, 2.0862e+05, -2.0715e+07, 1.3481e+07, 2.1496e+06, 5.6908e+06, 
    2.0731e+07, -1.7394e+07, 9.7651e+06, 6.0091e+06, -1.8077e+07, 
    -5.2843e+06, -5.139e+05, 5.4209e+06, -2.9637e+06, 8.7678e+05, 
    -2.3296e+07, 7.7239e+06, -7.6165e+06, 1.2251e+06, -3.0625e+06, 
    -3.0124e+06, 7.4043e+06, 3.5243e+06, -6.523e+06, 7.1347e+06, 9.0187e+06, 
    -7.8719e+06, -1.4852e+06, -1.3867e+07, 1.0832e+07, -1.8595e+06, 
    6.4704e+06, 2.2403e+06, 1.2587e+07, -3.5276e+06, -3.6175e+06, 2.8887e+07, 
    4.7071e+06, 4.5118e+06, -1.0409e+07, 1.1487e+07, 2.5752e+06,
  7.4408e+06, 3.3119e+06, -7.0537e+06, -3.0402e+07, -2.3156e+07, 4.3022e+06, 
    1.2709e+07, 3.3109e+07, -4.6254e+06, -9.5347e+06, 2.9282e+07, 2.0152e+07, 
    -3.1447e+07, -1.1502e+07, 3.4192e+05, 3.4007e+07, 2.6115e+07, 9.2736e+06, 
    -2.7133e+06, 1.5463e+07, 2.2115e+07, 2.5062e+07, 6.0843e+06, 1.0108e+07, 
    2.2417e+07, -5.7091e+06, 7.4937e+05, -2.6012e+07, 6.7669e+06, 3.1913e+07, 
    -1.9496e+05, 2.0102e+06, 2.5795e+07, -8.2978e+06, 8.203e+06, 3.0258e+06, 
    2.2988e+07, 1.5413e+07, -7.7016e+06, -7.9148e+06, 1.7023e+07, 3.4726e+06, 
    2.5975e+07, -1.6588e+07, 7.9902e+06, -2.1429e+07, 9.8224e+06, 
    -2.1484e+06, 2.8825e+06, -4.7607e+06, 1.7807e+07, 1.8551e+07, 
    -3.1132e+05, 7.0539e+06, -2.3266e+07, 1.5714e+06, 1.9073e+07, 
    -4.5156e+06, 16436, 3.0029e+07, -1.0129e+07, 1.8054e+07, 7.3062e+05, 
    1.3434e+07, -9.1588e+06, 1.6342e+06, -8.471e+06, -5.5321e+06, 
    -1.3263e+07, 6.2846e+06, 3.9383e+05, 1.7885e+07, -3.5812e+07, 7.8579e+06, 
    -6.6353e+06, -2.5554e+06, 2.5809e+07, 5.8137e+05, 9.2347e+05, 
    -3.8029e+06, 2.4356e+06, 5.5743e+06, 2.5193e+07, 9.8965e+05, -3.6896e+07, 
    -2.2611e+07, -2.7376e+06, 2.7085e+07, 1.2366e+06, -1.0622e+06, 
    -1.2516e+07, 1.1528e+07, -1.373e+07, -8.9678e+05, -2.4806e+07, 
    -1.0911e+06, -3.8932e+06, 1.8177e+07, 2.7586e+06, -8.1983e+06,
  -1.3883e+07, 2.4696e+07, -2.0472e+07, 1.1582e+07, -9.002e+06, 1.4298e+07, 
    1.7801e+07, 1.3774e+07, 1.4878e+07, -1.7203e+06, 1.417e+07, -2.1154e+07, 
    2.362e+07, -3.0132e+07, -2.6913e+07, 1.2209e+07, 2.3805e+07, 1.3416e+07, 
    3.0761e+06, 3.3052e+07, -2.8216e+07, 3.2295e+06, -1.1614e+07, 6.7665e+06, 
    1.6396e+07, 4.461e+06, 1.2769e+07, -5.0704e+06, -2.8618e+07, 2.5327e+07, 
    -2.1609e+07, -7.9995e+06, 1.0478e+07, 5.7167e+06, 2.4787e+07, 3.0309e+07, 
    1.1633e+07, -6.5136e+05, 1.5454e+07, 6.4491e+06, -1.6073e+07, 
    -8.6641e+06, -7.4741e+05, 2.4486e+07, -3.0394e+07, 2.3984e+07, 
    -2.3365e+07, 2.0826e+07, -9.134e+06, 2.633e+07, -1.7815e+06, -1.9474e+07, 
    -9.2893e+06, -9.5239e+06, -5.4627e+06, -1.8182e+07, 9.1405e+06, 
    -5.7971e+06, -1.134e+07, 1.1115e+07, -3.0089e+06, -1.9184e+07, 
    -1.037e+07, -3.2632e+07, -1.0344e+07, 5.7557e+06, -3.2017e+07, 
    -4.0703e+06, 1.9244e+07, 1.5978e+07, 4.4179e+06, 3.0917e+07, 2.1377e+07, 
    2.3838e+07, 2.2207e+07, -2.8843e+07, 5.1936e+06, 2.1998e+07, 4.1756e+07, 
    9.6915e+06, -1.4739e+07, -6.9238e+06, 1.1743e+07, -1.4469e+07, 
    -1.1973e+07, -1.7096e+07, 8.2229e+06, -5.2661e+06, -2.0241e+07, 
    2.3769e+07, 2.5793e+07, 8.7461e+06, 6.7791e+06, 5.8193e+06, 3.6266e+06, 
    -2.2021e+07, -2.3021e+07, 1.1934e+07, 2.8479e+07, 2.1652e+07 ;

 v_gns =
  4479.1, 1512.6, 51.809, -0.64232, -1682.8, 7660.5, -3992.5, 1685.9, 
    -1224.5, 382.6, -2350.2, -3575.6, -157.46, 2710.4, -2567, -962.14, 
    -1657.9, 228.29, 525.9, -2.7318, 3.4565, 1129.4, 2102.9, 1382.2, 224.8, 
    1563.1, 538.44, 365.46, 3242.9, 1477.9, 719.79, -2854.6, -156.99, 977.15, 
    306.59, 1111.2, 24.446, 5362.6, -5461.6, 1361.7, -4946.7, 2791, -612, 
    -3306.5, 17.802, 320.59, -1681.6, 761.25, 554.49, 205.61, -1039, 810.3, 
    -110.99, -1617.8, 2302.6, -1290.1, 8107.4, 232.59, -1306.8, 12.488, 
    694.08, 982.63, 339.14, 3563.1, 2793.3, 848.38, -5229.2, 3686.1, 289.07, 
    5811, -102.53, -4761.2, 2459.8, -5302.8, 4780, -3003.4, 781.92, -391.05, 
    -6373, 1735.1, -6480.4, 1198, -536.31, 914.56, 3528.4, -5949.4, 2160.1, 
    -364.46, -645.54, 5399.5, 742.96, 2921.9, -889.11, -522.36, 2563.9, 
    -4857, -277.29, 743.98, -1.5474, -901.91,
  -225.33, -1375.2, 1424.1, -12.466, 2102.3, 3642.6, 4010.8, -7963.6, 4595.5, 
    -1692.1, -1348.3, -2089.6, -3055.1, -2806.6, -580.95, 4045.4, 1622, 
    -176.02, -19.24, -0.21841, 76.236, 2622.4, -932.85, -180.21, -365.81, 
    3866.2, 4627, 288.72, 816, 1261.1, -278.54, -5138.4, 334.49, 1593.3, 
    633.24, -1189.1, -47.631, -7536.3, 1591.7, 6587.1, -2040.5, 5428.5, 
    580.45, -705.46, 21.579, -618.31, -4098.3, -2533.2, -116.31, 201.89, 
    1074.7, 796.35, -186.68, -3323.7, 615.51, -2028.1, -379.2, 4210.9, 
    4282.2, -2.3607, -41.77, -663.3, -1011.1, 3646.4, -1839.8, -134.26, 
    2720.3, -180.39, 537.99, 7117.4, -94.238, 3829.1, 1410.2, -2871.2, 
    -1461.8, -73.811, -532.8, -3337, -1887.4, 694.75, -3673.7, 2861.4, 
    836.82, 1860.4, 1053.3, 6341.1, 6889, 563.34, 6656, -3005, -2375.7, 
    2059.2, -2366, -8995.6, -8180.8, 1589.7, -429.5, 2407.8, 2.8965, 2506.7,
  -5418.8, -5423.2, -5589.3, -7172.7, -5880.1, -1179.5, 7694, 1156.9, 6749.6, 
    -5028.3, -5225.9, 5933.4, 179.25, -6681.7, 4688, -1836.1, -8634.6, 
    147.25, 182.05, -13.071, 111.75, 3174.2, 776.63, -1777.8, 49.988, 475.46, 
    6409.1, 1713.3, -2649.1, -4615, 3494.3, -4336, -411.69, 866.8, -1969.9, 
    3868.9, -146.46, 1530.3, 3134.4, -5819, 6.4148, 5684.4, -2584.3, 1502.7, 
    -9444.7, -2595.6, -4241.1, 3128.9, -3484, -6405.5, -6399.2, 338.53, 
    2223.3, -1901.5, -1952, -4653.4, -373.47, 771.12, 627.24, -1.3202, 
    345.24, -960.89, 6367, -6626.7, 112.44, -510.42, 1505, -5585.9, 1798.6, 
    -2430.8, -4087.7, 5794.9, -104.26, 3927.6, -2937.7, 523.37, -647.89, 
    -5490.2, -1999.6, -1671.4, -1127.8, 6571.8, 5326.8, -1102.9, -2814.5, 
    -2824.1, 6165.3, 8293.9, 1740.6, 23.554, 4909.5, 4881.9, 8569.3, -152.11, 
    -3398.2, -7640.2, -725.67, -3494.5, -8.3848, 3963.4 ;

 r_leo =
  -1.9449e+06, -3.3775e+06, 6.5888e+06, 6.5353e+06, -6.0101e+05, -3.5608e+06, 
    8.0953e+05, -4.9896e+06, 5.0645e+05, 3.2997e+06, -7.0392e+06, 1.1133e+05, 
    -2.151e+06, -1.3439e+06, 3.6443e+06, -2.1651e+06, 6.1654e+06, 5.2834e+06, 
    5.0008e+06, 8.2185e+05, 5.0136e+06, -55043, 4.0171e+06, 1.6935e+06, 
    6.2718e+06, 5.7534e+06, -3.7657e+06, 6.6094e+06, 6.5735e+05, -2.5866e+06, 
    6.823e+06, 4.4726e+06, -1.068e+05, 43493, -8.6112e+05, 3.9498e+06, 
    -41492, -2.8678e+05, 2.1234e+06, 1.5548e+06, -2.3498e+06, -4.9616e+06, 
    -4.4079e+06, -5.469e+06, 5.2178e+06, 5.2378e+06, -1.2475e+06, 
    -2.7369e+06, 3.4498e+06, -4.0072e+06, -6.4947e+06, 7.2184e+06, 
    -3.2804e+06, 5.076e+06, 8.6585e+06, -4.6216e+06, 4.318e+06, 1.435e+06, 
    2.4049e+06, 3.8077e+05, 2.5672e+06, -6.3264e+06, 9.5714e+05, -2.0235e+06, 
    -5.0788e+06, -8.9271e+05, 4.6151e+06, 1.2674e+06, 4.6383e+06, 1.1036e+06, 
    4.0104e+05, 5.1345e+06, -5.5199e+05, -3.3853e+06, 4.4666e+06, 
    -6.1954e+06, 1.0131e+05, -5.3334e+05, -2.5891e+06, -1.7803e+06, 
    6.265e+06, -5.0518e+06, -1.8793e+06, 3.5739e+06, 2.5585e+06, -6.99e+06, 
    -2.0018e+06, 2.4098e+06, 9.1707e+05, -2.0015e+06, 2.8716e+06, 1.6987e+06, 
    4.6494e+06, -3.0636e+06, 6.1562e+06, 2.2429e+06, -2.2958e+05, 
    -8.4331e+05, -7.492e+06, -90176,
  6.0482e+05, 9.2446e+05, -5.2353e+06, -5.6351e+06, -3.737e+06, 5.255e+06, 
    7.4145e+06, -6.0497e+06, -2.5152e+06, -5.5918e+06, 3.5265e+06, 
    2.3616e+05, 2.6836e+06, -2.0901e+06, 5.357e+06, -2.4736e+05, 1.1771e+06, 
    -3.5219e+06, 5.7122e+06, -6.8687e+06, -4.8166e+06, -7.1126e+05, 
    -1.8923e+06, 9.6471e+05, -1.3534e+06, -3.0718e+06, 1.497e+06, 
    -1.0032e+06, -6.3406e+06, 8.5323e+06, 4.026e+05, 5.7136e+06, 25969, 
    8.1076e+06, 5.9929e+06, 2.2618e+06, 7.1854e+05, 9.6545e+06, -1.3598e+06, 
    -6.1607e+06, 2.4328e+06, -5.5148e+06, -1.8422e+06, -5.1084e+06, 
    2.9246e+06, -5.6065e+06, 3.4349e+05, 1.7062e+06, -1.2643e+06, 
    -6.5515e+06, 2.7139e+06, -1.9608e+06, -3.3842e+06, -2.5141e+05, 
    5.8714e+05, -3.2315e+05, -5.7633e+06, -1.3745e+06, 1.0857e+06, 
    7.9597e+06, 1.8012e+06, 8.0653e+05, -7.5325e+06, -1.1387e+06, 2.6713e+06, 
    -8.0959e+05, -8.128e+05, 2.312e+06, 7.5106e+06, -8.657e+05, 9.2163e+06, 
    -4.1977e+06, 5.6004e+06, -2.3955e+06, -1.5419e+06, 1.6354e+06, 
    1.1062e+06, -5.9334e+06, -9.0892e+05, -3.2752e+06, -1.0123e+06, 
    -2.7646e+06, 6.1026e+06, 9.9062e+05, 1.9794e+06, -5.9251e+06, 
    -2.7902e+06, -2.6507e+06, 4.491e+06, -2.5416e+06, 4.3152e+06, 
    -2.4891e+06, 4.9234e+06, -1.8204e+06, -3.5313e+06, 8.4091e+06, 
    -3.9398e+05, -3.9093e+05, 2.3909e+06, -1.3847e+06,
  6.5616e+06, 6.7118e+06, 1.3912e+06, -4.4533e+06, -6.4233e+06, 1.1439e+06, 
    -6.4901e+06, -3.1644e+06, -5.8116e+06, -4.8452e+06, -2.3922e+06, 
    -9.2911e+06, 9.2491e+06, 8.4797e+06, -3.641e+06, 8.4502e+06, -2.0277e+06, 
    -4.8463e+06, 5.5782e+06, 3.0735e+06, -2.8377e+06, 8.3261e+06, 6.1287e+06, 
    7.1102e+06, -3.6508e+05, 1.7525e+05, -8.4066e+06, -7.1637e+06, 
    -6.0508e+05, -2.6504e+06, -2.2917e+06, -6.517e+06, -8.7792e+06, 
    -2.4686e+06, 5.7524e+06, -5.3802e+06, 8.7633e+06, -6.913e+05, 9.4019e+06, 
    5.0714e+06, -7.0531e+06, 3.5221e+06, -7.7717e+06, 2.7448e+06, 2.361e+06, 
    3.6971e+06, 6.366e+06, -8.6739e+06, 5.8149e+06, -2.0942e+06, 2.1216e+06, 
    -4.9034e+06, 4.7924e+06, 3.5563e+06, -4.3814e+06, -4.8963e+06, 
    -6.6619e+05, -5.9071e+06, -7.4631e+06, -1.2276e+05, 6.8942e+06, 
    -1.975e+06, 3.4925e+06, 9.1075e+06, 6.1023e+06, 7.1613e+06, -6.5425e+06, 
    -7.1099e+06, -4.4066e+06, 7.1507e+06, -8.2429e+05, -1.5203e+06, 
    -5.2015e+06, 5.1542e+06, -8.1067e+06, -6.8338e+06, 7.5001e+06, 
    -6.738e+06, -5.8769e+06, -5.9758e+06, -6.4009e+06, 4.4645e+06, 
    4.9191e+06, 8.7773e+06, -5.4089e+06, 1.9651e+06, 9.2171e+06, 6.2593e+06, 
    -7.0557e+06, 5.3782e+06, 3.749e+06, -6.4362e+06, -4.1349e+06, 7.4171e+06, 
    6.2968e+06, -2.65e+06, -9.5416e+06, -6.2091e+06, 1.273e+06, 8.6481e+06 ;

 v_leo =
  1333, 543.16, 474.68, 3343.9, -309.38, -38.94, 5132.1, 3653, -7322.9, 
    4618.7, 2896, -634.54, 3170.6, -288.94, -9.6591, -3472.8, -5008, 900.91, 
    -5593.4, 6893.4, 509.4, 3037.8, -892.82, 1944.2, 2986.3, 3421.9, -3570.7, 
    -248.34, -453.6, -2152.5, -2.7605, 390.21, -3337.6, 4718.6, -3777.5, 
    8836.4, 623.4, 1266.4, -592.57, -876.38, 547.7, 728.78, -588.72, -4668.5, 
    -56.408, -3710.4, -194.26, -938.07, -562.25, -8003.5, 2061.2, 1121.1, 
    878.17, -708.62, -1546.1, -68.379, -3677.9, -357.14, 3.2423, -319.85, 
    -2801.3, -1131.5, 484.81, -1415.2, -198.87, -2872.6, -652.88, -195.27, 
    -3999.7, 2266, 1333.8, -2466, 4536.2, -1056.3, 6753, -89.561, -2182.2, 
    -810.39, 241.71, 6610.5, -518.91, 976.47, -5003.3, -1060.9, 509.49, 
    -1572.9, -441.06, -3104, 89.881, 4726.5, -472.39, 6053.4, 2849.2, 
    -942.89, -3455.2, -673.87, 704.65, -3303.8, 8631.5, 2939.1,
  721.28, -81.061, -340.77, -3272.5, -2483.5, -1793.6, 2318.1, -126.74, 
    -3159, 667.56, -3804.9, 2890, -4332, 629.95, 34.621, 483.41, -3301.8, 
    -6751.9, -2585.5, 3005.4, -2322.5, -823.19, -470.35, 4185.4, 4539.7, 
    4080.8, -7119.2, -4267.3, -278.09, -3687.9, 14.408, 176.35, -2704.8, 
    -3570.1, 4708.4, 1620.5, 5352.7, 3721.4, -5209, 1296.3, -3158.2, 1227.3, 
    -2467.5, 4493.4, 614.73, -5226.2, -2787.6, 306.92, -2722.5, 3031.7, 
    2199.7, -718.49, -527.67, -1125, -1767.1, 463.15, -3449.2, 688.86, 58.6, 
    2743.3, 3142.1, 1406.9, -1530.4, -1381.8, -805.65, -6001.1, -600.5, 
    609.34, -1999.5, 5518.9, -7042.6, 4776.5, -1582.2, 583.21, -4461.6, 
    -106.75, 3441.8, 379.08, -1426, 3594.1, 685.26, 112.45, 746.12, -1429.5, 
    -2478, 1253.7, -477.02, 1957.1, 46.436, -7791.4, -6533.7, 376.21, 2713.2, 
    -309.07, -3575.4, -111.9, 273.2, -450.49, 987.13, 6454.1,
  885.73, 7592.4, -1128.6, -3983.8, -2901.1, 7866.8, 5719.2, 5008.8, -3595.1, 
    -982.06, 4295.1, 1049.7, -4537.7, -1036.5, 24.456, 4919.8, 4041.3, 
    1964.2, -1196.4, 2818.5, 1045.9, 4372, 1179, 5090.1, 4372.6, -4694, 
    316.01, -1656.5, 513.62, 5642.5, -69.804, 901.15, 4507.6, -2885.4, 
    6646.2, 3024.8, 3378.7, 2877.9, -6679.3, -6004.3, 1054, 642.17, 4214.5, 
    -4749.4, 546.05, -3862.9, 489.09, -8585.3, 368.25, -2089.7, 3589.4, 
    2283.8, -51.545, 1558.1, -3636.9, 142.66, 3914.8, -3226, 2.3082, 5260.4, 
    -1405.2, 1603.3, 102.63, 584.83, -3357.1, 552.86, -458.32, -4277.4, 
    -6595.2, 6473.8, 260.03, 6339.6, -4688.1, 7352.6, -2999.1, -853.39, 
    3886.5, 9509.9, 9652.5, -1819.3, 268.12, 2663.2, 3825, 97.376, -3126.5, 
    -2147.8, -6645.5, 2484.5, 334.82, -743.02, -5482.3, 2357.8, -5073, 
    -8126.4, -1841.9, -78.136, -281, 5751.9, 1028.6, -5205.8 ;

 phase_qual =
  27.445, 74.881, 43.533, 72.559, 51.304, 30.445, 42.589, 84.769, 26.923, 
    47.609, 71.964, 87.336, 90.996, 71.744, 56.291, 86.39, 83.391, 42.894, 
    4.5558, 93.397, 95.069, 55.502, 18.873, 16.315, 59.794, 2.9382, 26.333, 
    88.948, 63.066, 96.539, 41.887, 6.0034, 58.884, 15.714, 54.134, 66.627, 
    59.411, 27.125, 30.35, 30.577, 72.502, 9.8603, 63.052, 64.77, 68.594, 
    75.804, 84.181, 45.317, 22.153, 60.009, 32.517, 61.61, 9.7649, 15.502, 
    54.094, 33.15, 42.135, 14.397, 13.973, 86.784, 29.696, 54.976, 15.357, 
    94.369, 43.514, 14.273, 74.619, 35.7, 48.264, 29.83, 2.1854, 80.543, 
    96.513, 76.209, 49.539, 64.512, 54.768, 43.527, 96.943, 17.868, 24.86, 
    13.113, 61.132, 29.561, 90.71, 60.287, 27.589, 63.701, 38.488, 50.153, 
    61.294, 35.269, 25.852, 1.9307, 87.088, 44.415, 47.77, 48.661, 66.934, 
    46.452 ;

 lat_tp =
  -18.295, -12.508, 77.794, -74.461, -38.202, 86.114, -66.407, 51.139, 
    -36.335, 57.063, -2.6971, 59.425, -68.584, -53.323, 28.365, -80.037, 
    59.001, -85.074, -20.052, 23.846, 61.312, 70.805, 13.29, -72.197, 6.1712, 
    -5.087, 2.6324, -18.949, 9.8207, -69.078, -53.247, -89.33, -73.733, 
    -77.988, -84.997, -61.162, 35.987, -4.5032, 67.005, -53.473, 82.773, 
    -53.968, -16.033, -66.86, 67.157, -48.504, -63.204, -73.24, 66.197, 
    -49.322, 58.636, -3.1396, 68.009, -70.417, -13.588, 0.45203, -71.652, 
    -34.376, -71.574, -39.166, -67.775, 49.258, -21.658, -82.245, 27.768, 
    23.146, 67.906, -12.262, 34.786, 55.136, -6.0936, -32.328, 74.218, 
    63.574, -9.8117, -52.91, 72.178, 34.705, -28.617, -25.372, 45.208, 
    -50.878, -40.951, 78.2, -27.752, 41.744, 37.866, 30.108, -36.107, 19.608, 
    -68.15, -10.061, -33.428, -85.133, -21.275, -49.336, 85.195, 66.012, 
    -70.46, -34.67 ;

 lon_tp =
  58.291, 65.462, 65.729, -44.605, -82.59, -55.904, -96.678, -107.91, 17.313, 
    -161.38, -10.92, 65.873, 69.739, 169.78, -33.474, 156.6, -53.469, 
    -128.39, -39.351, 119.18, 120.32, -112.69, 44.713, 131.32, -47.956, 
    76.547, -4.5725, 21.837, -15.682, 10.094, 33.739, 159.5, 118.02, -51.172, 
    121.73, 3.2407, -132.08, -139.88, -116.77, 89.976, -26.063, 30.939, 
    -104.53, 55.33, -54.518, 65.048, -165.29, -11.637, -30.644, -66.7, 72.66, 
    108.39, -169.3, 155.35, 119.77, -102.59, -60.602, -170.7, 55.922, 49.81, 
    10.371, 0.16601, -144.45, 70.144, -65.825, -139.78, -68.697, -89.036, 
    3.4661, 120.69, 76.759, 49.542, 106.57, 33.241, -95.561, 162.65, 91.202, 
    15.012, 108.5, 4.632, -13.402, 163.08, 148.2, -92.993, -174.09, -48.38, 
    -13.432, 45.412, -12.732, 98.243, -48.354, -93.087, -132.24, 57.81, 
    -34.323, 69.067, 121.24, 105.13, 80.175, 126.99 ;

 azimuth_tp =
  186.34, 18.795, 316.01, 301.69, 12.03, 110.11, 107.33, 219.07, 36.365, 
    98.089, 47.515, 351.84, 212.16, 133.95, 21.405, 111.37, 195.01, 250.78, 
    307.8, 81.362, 239.88, 58.594, 56.714, 348.14, 73.858, 340.11, 40.681, 
    63.664, 137.59, 351.58, 85.824, 118.05, 52.017, 203.7, 1.1575, 318.46, 
    60.073, 109.88, 79.659, 101.23, 78.557, 130.79, 178.35, 6.5388, 128.04, 
    38.754, 319.02, 328.56, 152.66, 322.73, 131.38, 110.99, 191.24, 59.479, 
    259.3, 178.73, 307.41, 25.217, 300.4, 167.29, 47.871, 58.547, 111.75, 
    185.46, 227.18, 259.17, 266.77, 315.09, 296.76, 186.25, 268.18, 120.23, 
    98.381, 254.19, 3.8721, 275.36, 89.258, 210.69, 182.1, 196.91, 332.39, 
    154.29, 311.58, 258.4, 277.86, 139.96, 175.53, 250.97, 161.04, 243.12, 
    6.0223, 205.16, 326.33, 7.4282, 150.18, 15.464, 192.96, 300.38, 230.3, 
    309.6 ;

 impact_L1 =
  6.5222e+06, 6.2529e+06, 6.5382e+06, 6.497e+06, 6.3905e+06, 6.4026e+06, 
    6.5523e+06, 6.3058e+06, 6.4947e+06, 6.2461e+06, 6.2892e+06, 6.2381e+06, 
    6.4166e+06, 6.4265e+06, 6.2476e+06, 6.2389e+06, 6.3149e+06, 6.3896e+06, 
    6.5764e+06, 6.5336e+06, 6.2305e+06, 6.2883e+06, 6.4686e+06, 6.5517e+06, 
    6.4975e+06, 6.5388e+06, 6.3886e+06, 6.2518e+06, 6.5799e+06, 6.2198e+06, 
    6.2091e+06, 6.2376e+06, 6.5623e+06, 6.4322e+06, 6.2125e+06, 6.4154e+06, 
    6.2628e+06, 6.3133e+06, 6.3457e+06, 6.373e+06, 6.3116e+06, 6.4896e+06, 
    6.4127e+06, 6.5784e+06, 6.4473e+06, 6.4601e+06, 6.2847e+06, 6.2222e+06, 
    6.3032e+06, 6.333e+06, 6.3908e+06, 6.5866e+06, 6.4177e+06, 6.4157e+06, 
    6.4976e+06, 6.4247e+06, 6.2343e+06, 6.4785e+06, 6.2999e+06, 6.5592e+06, 
    6.3085e+06, 6.3145e+06, 6.3424e+06, 6.214e+06, 6.4874e+06, 6.3509e+06, 
    6.4141e+06, 6.5571e+06, 6.3093e+06, 6.2848e+06, 6.3985e+06, 6.5581e+06, 
    6.2314e+06, 6.4296e+06, 6.2405e+06, 6.3871e+06, 6.4971e+06, 6.3843e+06, 
    6.4498e+06, 6.5878e+06, 6.3174e+06, 6.2331e+06, 6.2455e+06, 6.3821e+06, 
    6.4866e+06, 6.535e+06, 6.4494e+06, 6.536e+06, 6.3573e+06, 6.5169e+06, 
    6.5064e+06, 6.5571e+06, 6.3068e+06, 6.5184e+06, 6.2269e+06, 6.515e+06, 
    6.2653e+06, 6.5521e+06, 6.2943e+06, 6.4056e+06 ;

 impact_L2 =
  6.5399e+06, 6.5047e+06, 6.2888e+06, 6.4705e+06, 6.4759e+06, 6.5044e+06, 
    6.434e+06, 6.2332e+06, 6.2252e+06, 6.2908e+06, 6.4107e+06, 6.2952e+06, 
    6.4991e+06, 6.2892e+06, 6.3523e+06, 6.4799e+06, 6.5395e+06, 6.4629e+06, 
    6.4531e+06, 6.2392e+06, 6.5881e+06, 6.497e+06, 6.565e+06, 6.339e+06, 
    6.5012e+06, 6.5679e+06, 6.4045e+06, 6.2969e+06, 6.2957e+06, 6.5687e+06, 
    6.4188e+06, 6.5686e+06, 6.5779e+06, 6.5099e+06, 6.2212e+06, 6.375e+06, 
    6.4952e+06, 6.2538e+06, 6.4599e+06, 6.4496e+06, 6.578e+06, 6.215e+06, 
    6.4669e+06, 6.5358e+06, 6.2237e+06, 6.2664e+06, 6.2894e+06, 6.275e+06, 
    6.2836e+06, 6.3939e+06, 6.3279e+06, 6.519e+06, 6.4539e+06, 6.4845e+06, 
    6.5086e+06, 6.2762e+06, 6.2384e+06, 6.5234e+06, 6.2389e+06, 6.4915e+06, 
    6.5257e+06, 6.5032e+06, 6.4966e+06, 6.4007e+06, 6.3901e+06, 6.524e+06, 
    6.4913e+06, 6.5176e+06, 6.258e+06, 6.5567e+06, 6.4048e+06, 6.4268e+06, 
    6.5377e+06, 6.3392e+06, 6.5498e+06, 6.4397e+06, 6.3548e+06, 6.3053e+06, 
    6.3908e+06, 6.4099e+06, 6.5677e+06, 6.3356e+06, 6.2218e+06, 6.4201e+06, 
    6.2412e+06, 6.3462e+06, 6.3837e+06, 6.5175e+06, 6.5735e+06, 6.3853e+06, 
    6.5747e+06, 6.2616e+06, 6.3075e+06, 6.3703e+06, 6.4353e+06, 6.3605e+06, 
    6.3502e+06, 6.4173e+06, 6.3383e+06, 6.5464e+06 ;

 impact =
  6.224e+06, 6.2569e+06, 6.2553e+06, 6.3537e+06, 6.5336e+06, 6.2863e+06, 
    6.3885e+06, 6.5495e+06, 6.5044e+06, 6.5711e+06, 6.4367e+06, 6.2037e+06, 
    6.4551e+06, 6.2426e+06, 6.3311e+06, 6.5852e+06, 6.3028e+06, 6.4895e+06, 
    6.2021e+06, 6.4417e+06, 6.5144e+06, 6.5311e+06, 6.5558e+06, 6.5234e+06, 
    6.5759e+06, 6.505e+06, 6.4653e+06, 6.3765e+06, 6.2284e+06, 6.3817e+06, 
    6.387e+06, 6.2538e+06, 6.4149e+06, 6.2211e+06, 6.4339e+06, 6.4854e+06, 
    6.3271e+06, 6.3502e+06, 6.5855e+06, 6.2054e+06, 6.2949e+06, 6.2083e+06, 
    6.4448e+06, 6.2978e+06, 6.3998e+06, 6.3173e+06, 6.5546e+06, 6.3895e+06, 
    6.3498e+06, 6.2239e+06, 6.5554e+06, 6.427e+06, 6.4122e+06, 6.562e+06, 
    6.231e+06, 6.3005e+06, 6.5408e+06, 6.5605e+06, 6.2383e+06, 6.2261e+06, 
    6.571e+06, 6.2978e+06, 6.5464e+06, 6.5438e+06, 6.4995e+06, 6.3231e+06, 
    6.2996e+06, 6.2534e+06, 6.4183e+06, 6.5802e+06, 6.3626e+06, 6.4825e+06, 
    6.5444e+06, 6.3633e+06, 6.51e+06, 6.5375e+06, 6.4675e+06, 6.566e+06, 
    6.4334e+06, 6.3912e+06, 6.3433e+06, 6.3444e+06, 6.5504e+06, 6.2582e+06, 
    6.4295e+06, 6.5552e+06, 6.4326e+06, 6.4723e+06, 6.2223e+06, 6.4148e+06, 
    6.512e+06, 6.2991e+06, 6.4987e+06, 6.4465e+06, 6.2404e+06, 6.4733e+06, 
    6.3026e+06, 6.3679e+06, 6.4372e+06, 6.3599e+06 ;

 impact_opt =
  6.3526e+06, 6.3285e+06, 6.4421e+06, 6.3729e+06, 6.5338e+06, 6.5261e+06, 
    6.5671e+06, 6.4019e+06, 6.3164e+06, 6.3194e+06, 6.3148e+06, 6.4179e+06, 
    6.5751e+06, 6.3561e+06, 6.3079e+06, 6.419e+06, 6.3553e+06, 6.4724e+06, 
    6.3458e+06, 6.3561e+06, 6.5581e+06, 6.2228e+06, 6.4122e+06, 6.5468e+06, 
    6.2659e+06, 6.263e+06, 6.3738e+06, 6.5248e+06, 6.3509e+06, 6.3188e+06, 
    6.2784e+06, 6.5418e+06, 6.2027e+06, 6.3496e+06, 6.3766e+06, 6.5073e+06, 
    6.4047e+06, 6.2535e+06, 6.5903e+06, 6.2302e+06, 6.3265e+06, 6.4586e+06, 
    6.4641e+06, 6.2019e+06, 6.4334e+06, 6.3844e+06, 6.5438e+06, 6.3039e+06, 
    6.2101e+06, 6.2658e+06, 6.4541e+06, 6.2912e+06, 6.456e+06, 6.5576e+06, 
    6.2025e+06, 6.5153e+06, 6.5675e+06, 6.2105e+06, 6.5222e+06, 6.3761e+06, 
    6.2081e+06, 6.3969e+06, 6.4142e+06, 6.4512e+06, 6.4228e+06, 6.2835e+06, 
    6.3835e+06, 6.4461e+06, 6.3188e+06, 6.4271e+06, 6.4165e+06, 6.2783e+06, 
    6.4698e+06, 6.4413e+06, 6.5388e+06, 6.5184e+06, 6.3277e+06, 6.2111e+06, 
    6.5612e+06, 6.4773e+06, 6.4223e+06, 6.5646e+06, 6.3336e+06, 6.507e+06, 
    6.2627e+06, 6.4734e+06, 6.2986e+06, 6.4218e+06, 6.4702e+06, 6.4436e+06, 
    6.5248e+06, 6.2621e+06, 6.2985e+06, 6.2737e+06, 6.5057e+06, 6.2975e+06, 
    6.3155e+06, 6.3823e+06, 6.2707e+06, 6.4802e+06 ;

 bangle_L1 =
  0.013973, 0.081249, 0.059904, 0.029306, 0.010693, 0.08019, 0.081691, 
    0.0084833, 0.04644, 0.081025, 0.0030973, 0.086541, 0.015102, 0.086824, 
    0.030157, 0.0029417, 0.023653, 0.0085311, 0.082219, 0.067257, 0.087362, 
    0.011568, 0.044546, 0.04711, 0.040502, 0.061493, 0.021367, 0.052821, 
    0.028934, 0.052338, 0.084815, 0.06988, 0.068877, 0.074664, 0.082024, 
    0.012381, 0.082073, 0.010393, 0.093103, 0.07321, 0.090365, 0.090506, 
    -0.00047212, 0.087305, 0.0072592, 0.027179, 0.041516, 0.097326, 0.078855, 
    0.063711, 0.0011314, 0.0075473, 0.067948, 0.092915, 0.050456, 0.069141, 
    0.0062308, 0.023423, 0.066425, 0.057174, 0.0019803, 0.075536, 
    -0.00095218, 0.040883, 0.07612, 0.061155, 0.093178, 0.024905, 0.044494, 
    0.024049, 0.049789, 0.07977, 0.059142, 0.093555, 0.040615, 0.020458, 
    0.042848, -0.00053665, 0.041949, 0.019352, 0.084609, 0.022863, 0.048105, 
    0.044284, 0.08261, 0.056595, 0.040997, 0.050706, 0.071496, 0.052629, 
    0.071914, 0.060335, 0.014811, 0.080933, 0.018888, 0.079811, 0.057181, 
    0.050588, 0.080274, 0.064211 ;

 bangle_L2 =
  0.0022921, 0.0066008, 0.065718, 0.088792, 0.074647, 0.076138, 0.096031, 
    0.013045, -0.00085846, 0.026525, 0.017181, 0.095314, 0.057047, 0.084814, 
    0.083403, 0.09194, 0.012745, 0.084369, 0.058254, 0.086232, 0.044866, 
    0.04498, 0.0077488, 0.030305, 0.0088659, 0.031201, 0.081406, 0.096658, 
    0.065379, 0.054573, 0.00020353, 0.017876, 0.079928, 0.0083745, 
    -0.00013444, 0.022548, 0.070829, 0.033415, 0.039176, 0.012045, 0.063404, 
    0.064631, 0.046866, 0.059381, 0.068837, 0.055147, 0.077527, 0.058849, 
    0.068685, 0.047086, 0.080594, 0.057738, 0.055376, 0.013848, 0.087704, 
    0.016484, 0.055402, 0.052214, 0.029336, 0.085514, 0.080677, 0.052067, 
    0.016351, 0.085506, 0.065907, 0.07564, 0.028302, 0.04076, 0.0074748, 
    0.047445, 0.035273, 0.031696, 0.038887, 0.024165, 0.034081, 0.036205, 
    0.018715, 0.051758, 0.042597, 0.072889, 0.065595, 0.096699, 0.071363, 
    0.071127, 0.078135, 0.073052, 0.046153, 0.061108, 0.085059, 0.083277, 
    0.001432, 0.046155, 0.089954, 0.017665, 0.009736, 0.062573, 0.017001, 
    0.052409, 0.014335, 0.066698 ;

 bangle =
  0.042304, 0.074392, 0.083104, 0.081512, 0.036908, 0.060801, 0.051545, 
    0.051081, 0.023452, 0.046876, 0.040812, 0.075272, 0.020246, 0.093545, 
    0.045187, 0.0059381, 0.056214, 0.033543, 0.046069, 0.028556, 0.048778, 
    0.011452, 0.0098735, 0.017668, 0.012798, 0.0372, 0.094801, 0.011211, 
    0.040254, 0.066259, 0.029034, 0.067519, 0.036335, 0.097215, 0.0022357, 
    0.087189, 0.019466, 0.078053, 0.084065, 0.032983, 0.044673, 0.079723, 
    0.085074, 0.046045, 0.080696, -0.00026308, 0.018595, 0.07576, 0.028713, 
    0.042581, 0.083506, 0.09709, 0.084399, 0.029095, 0.00031572, 0.095698, 
    0.018251, 0.076794, 0.096349, 0.093657, 0.0088767, 0.061286, 0.080452, 
    0.085556, 0.074689, 0.069137, 0.010083, 0.0090962, 0.061456, 0.00030602, 
    0.081974, 0.0034517, 0.022764, 0.011615, 0.015409, -0.0001736, 0.089451, 
    0.076637, 0.084547, 0.021925, 0.034633, 0.02008, 0.075392, 0.033145, 
    0.087744, 0.096486, 0.088888, 0.0017462, 0.093047, 0.041628, 0.079865, 
    0.089042, 0.072617, 0.043513, 0.028559, 0.029768, 0.050955, 0.031819, 
    0.046165, 0.09625 ;

 bangle_opt =
  0.039234, 0.042482, 0.093151, 0.0077189, 0.028064, 0.097819, 0.012238, 
    0.078195, 0.029112, 0.081519, 0.047987, 0.082844, 0.011017, 0.01958, 
    0.065416, 0.0045901, 0.082606, 0.001764, 0.038248, 0.06288, 0.083903, 
    0.089229, 0.056957, 0.0089897, 0.052963, 0.046646, 0.050977, 0.038867, 
    0.055011, 0.010739, 0.019622, -0.0006238, 0.0081276, 0.0057401, 0.001807, 
    0.015181, 0.069693, 0.046973, 0.087097, 0.019496, 0.095945, 0.019218, 
    0.040504, 0.011984, 0.087183, 0.022284, 0.014036, 0.0084044, 0.086644, 
    0.021825, 0.082401, 0.047738, 0.087661, 0.0099881, 0.041876, 0.049754, 
    0.0092951, 0.030211, 0.009339, 0.027523, 0.011471, 0.077139, 0.037347, 
    0.0033517, 0.065081, 0.062487, 0.087603, 0.04262, 0.069019, 0.080437, 
    0.046081, 0.03136, 0.091145, 0.085172, 0.043995, 0.019812, 0.09, 
    0.068974, 0.033442, 0.035263, 0.074867, 0.020952, 0.026522, 0.093379, 
    0.033928, 0.072923, 0.070747, 0.066394, 0.02924, 0.060503, 0.01126, 
    0.043855, 0.030743, 0.0017309, 0.037562, 0.021817, 0.097304, 0.08654, 
    0.0099641, 0.030046 ;

 bangle_L1_sigma =
  0.0062783, 0.0064673, 0.0064743, 0.0035673, 0.0025665, 0.0032696, 
    0.0021953, 0.0018992, 0.0051986, 0.00049047, 0.0044548, 0.0064781, 
    0.0065799, 0.0092157, 0.0038606, 0.0088684, 0.0033338, 0.0013598, 
    0.0037057, 0.0078826, 0.0079126, 0.0017735, 0.0059206, 0.0082024, 
    0.003479, 0.0067593, 0.004622, 0.0053178, 0.0043293, 0.0050084, 
    0.0056314, 0.0089449, 0.007852, 0.0033943, 0.0079498, 0.0048279, 
    0.0012626, 0.0010569, 0.001666, 0.0071131, 0.0040558, 0.0055577, 
    0.0019885, 0.0062003, 0.0033061, 0.0064563, 0.00038762, 0.0044359, 
    0.0039351, 0.0029851, 0.0066569, 0.0075983, 0.00028204, 0.0088356, 
    0.0078982, 0.0020395, 0.0031458, 0.00024497, 0.0062159, 0.0060548, 
    0.0050158, 0.0047469, 0.00093655, 0.0065906, 0.0030082, 0.0010596, 
    0.0029325, 0.0023966, 0.0048338, 0.0079224, 0.0067649, 0.0060478, 
    0.0075502, 0.0056183, 0.0022247, 0.0090278, 0.0071454, 0.005138, 
    0.0076011, 0.0048645, 0.0043894, 0.0090393, 0.0086473, 0.0022924, 
    0.00015571, 0.0034678, 0.0043886, 0.005939, 0.004407, 0.0073309, 
    0.0034685, 0.0022899, 0.0012583, 0.0062656, 0.0038382, 0.0065622, 
    0.0079368, 0.0075124, 0.0068549, 0.0080883 ;

 bangle_L2_sigma =
  0.0049095, 0.00049518, 0.0083259, 0.0079486, 0.00031695, 0.002901, 
    0.0028278, 0.0057719, 0.00095813, 0.0025844, 0.0012519, 0.0092699, 
    0.0055898, 0.0035293, 0.00056396, 0.0029344, 0.0051379, 0.0066073, 
    0.0081096, 0.0021437, 0.0063201, 0.0015438, 0.0014943, 0.0091726, 
    0.001946, 0.0089609, 0.0010718, 0.0016774, 0.0036251, 0.0092631, 
    0.0022612, 0.0031102, 0.0013705, 0.0053668, 3.0496e-05, 0.0083905, 
    0.0015828, 0.0028951, 0.0020988, 0.0026672, 0.0020698, 0.0034458, 
    0.004699, 0.00017228, 0.0033736, 0.0010211, 0.0084054, 0.0086567, 
    0.0040221, 0.0085031, 0.0034614, 0.0029242, 0.0050385, 0.0015671, 
    0.0068318, 0.004709, 0.0080995, 0.00066439, 0.0079147, 0.0044077, 
    0.0012613, 0.0015425, 0.0029442, 0.0048863, 0.0059856, 0.0068285, 
    0.0070287, 0.0083017, 0.0078188, 0.0049073, 0.0070658, 0.0031678, 
    0.0025921, 0.0066972, 0.00010202, 0.007255, 0.0023517, 0.0055511, 
    0.0047979, 0.0051881, 0.0087575, 0.004065, 0.0082094, 0.0068082, 
    0.007321, 0.0036874, 0.0046246, 0.0066124, 0.0042428, 0.0064056, 
    0.00015867, 0.0054053, 0.0085978, 0.00019571, 0.0039569, 0.00040743, 
    0.0050838, 0.0079142, 0.0060678, 0.0081571 ;

 bangle_sigma =
  0.0076408, 0.0012549, 0.0080187, 0.0070435, 0.0045167, 0.0048051, 0.008355, 
    0.0025084, 0.0069875, 0.001094, 0.002116, 0.00090227, 0.005136, 0.005372, 
    0.0011284, 0.00092169, 0.0027247, 0.0044951, 0.0089246, 0.0079102, 
    0.00072346, 0.0020948, 0.0063682, 0.0083403, 0.0070556, 0.0080338, 
    0.0044717, 0.001228, 0.0090093, 0.00046965, 0.00021637, 0.00089173, 
    0.0085902, 0.005507, 0.00029654, 0.0051087, 0.0014893, 0.002687, 
    0.0034544, 0.0041022, 0.0026468, 0.0068668, 0.0050443, 0.0089727, 
    0.0058647, 0.0061668, 0.0020093, 0.00052724, 0.0024478, 0.0031545, 
    0.0045252, 0.0091675, 0.005163, 0.0051153, 0.0070563, 0.0053275, 
    0.00081434, 0.0066045, 0.0023685, 0.0085168, 0.0025724, 0.0027146, 
    0.0033761, 0.00033237, 0.0068154, 0.0035791, 0.0050777, 0.0084666, 
    0.0025906, 0.0020109, 0.0047058, 0.0084908, 0.00074458, 0.0054435, 
    0.00096017, 0.0044377, 0.0070443, 0.00437, 0.0059232, 0.0091958, 
    0.0027848, 0.00078415, 0.0010791, 0.0043183, 0.0067957, 0.0079448, 
    0.0059146, 0.0079679, 0.0037298, 0.0075146, 0.0072663, 0.0084672, 
    0.0025323, 0.0075494, 0.00063788, 0.007469, 0.0015478, 0.0083482, 
    0.0022369, 0.0048746 ;

 bangle_opt_sigma =
  0.0084973, 0.0076177, 0.0022189, 0.0067619, 0.0068977, 0.0076089, 
    0.0058509, 0.0008308, 0.00062881, 0.0022689, 0.0052672, 0.002379, 
    0.0074781, 0.0022294, 0.0038067, 0.0069966, 0.0084879, 0.0065736, 
    0.0063275, 0.00098095, 0.0097026, 0.0074245, 0.0091252, 0.0034754, 
    0.0075303, 0.0091963, 0.0051133, 0.0024218, 0.0023915, 0.0092165, 
    0.0054694, 0.0092155, 0.0094481, 0.0077475, 0.00052923, 0.0043759, 
    0.0073812, 0.0013442, 0.0064983, 0.0062391, 0.0094509, 0.00037493, 
    0.0066713, 0.0083956, 0.00059369, 0.0016599, 0.0022357, 0.0018738, 
    0.0020896, 0.0048466, 0.0031982, 0.0079753, 0.0063482, 0.0071129, 
    0.007716, 0.0019044, 0.00095902, 0.0080862, 0.00097303, 0.0072878, 
    0.0081425, 0.0075796, 0.0074142, 0.0050167, 0.0047533, 0.0080998, 
    0.0072834, 0.0079401, 0.001451, 0.0089167, 0.0051199, 0.0056702, 
    0.0084437, 0.0034808, 0.0087456, 0.0059933, 0.0038691, 0.0026322, 
    0.0047694, 0.0052486, 0.0091924, 0.0033909, 0.00054574, 0.0055027, 
    0.0010298, 0.0036548, 0.0045934, 0.0079369, 0.009337, 0.0046328, 
    0.0093676, 0.0015405, 0.0026881, 0.0042583, 0.0058833, 0.0040127, 
    0.0037554, 0.005432, 0.0034576, 0.0086606 ;

 bangle_L1_qual =
  5.9979, 14.236, 13.815, 38.415, 83.405, 21.572, 47.116, 87.376, 76.098, 
    92.775, 59.18, 0.93659, 63.77, 10.643, 32.777, 96.312, 25.702, 72.366, 
    0.51812, 60.431, 78.6, 82.764, 88.948, 80.846, 93.981, 76.244, 66.333, 
    44.121, 7.1118, 45.421, 46.751, 13.454, 53.734, 5.2717, 58.48, 71.347, 
    31.772, 37.557, 96.371, 1.361, 23.726, 2.0804, 61.193, 24.44, 49.947, 
    29.323, 88.658, 47.386, 37.441, 5.9648, 88.841, 56.756, 53.05, 90.503, 
    7.7394, 25.113, 85.202, 90.135, 9.587, 6.5145, 92.757, 24.44, 86.599, 
    85.943, 74.871, 30.779, 24.91, 13.349, 54.57, 95.062, 40.655, 70.624, 
    86.105, 40.816, 77.506, 84.384, 66.878, 91.502, 58.356, 47.804, 35.828, 
    36.101, 87.606, 14.552, 57.37, 88.804, 58.145, 68.077, 5.5634, 53.71, 
    78.007, 24.781, 74.667, 61.635, 10.104, 68.323, 25.653, 41.973, 59.295, 
    39.985 ;

 bangle_L2_qual =
  38.147, 32.127, 60.532, 43.224, 83.456, 81.521, 91.772, 50.469, 29.111, 
    29.838, 28.708, 54.484, 93.787, 39.024, 26.969, 54.748, 38.824, 68.094, 
    36.456, 39.03, 89.514, 5.7095, 53.046, 86.688, 16.467, 15.745, 43.447, 
    81.193, 37.733, 29.691, 19.592, 85.446, 0.67324, 37.396, 44.139, 76.816, 
    51.176, 13.383, 97.573, 7.557, 31.635, 64.648, 66.027, 0.46841, 58.346, 
    46.1, 85.939, 25.982, 2.5147, 16.453, 63.52, 22.795, 63.995, 89.404, 
    0.61321, 78.825, 91.873, 2.637, 80.543, 44.036, 2.0308, 49.236, 53.546, 
    62.804, 55.701, 20.885, 45.884, 61.526, 29.711, 56.777, 54.129, 19.583, 
    67.446, 60.329, 84.711, 79.605, 31.916, 2.7693, 90.308, 69.334, 55.574, 
    91.161, 33.392, 76.76, 15.678, 68.34, 24.656, 55.462, 67.562, 60.9, 
    81.209, 15.523, 24.63, 18.415, 76.434, 24.374, 28.885, 45.577, 17.682, 
    70.06 ;

 bangle_qual =
  14.825, 81.434, 60.301, 30.006, 11.577, 80.386, 81.872, 9.3894, 46.97, 
    81.212, 4.0567, 86.674, 15.943, 86.955, 30.848, 3.9027, 24.408, 9.4367, 
    82.395, 67.581, 87.487, 12.444, 45.095, 47.634, 41.091, 61.875, 22.145, 
    53.288, 29.637, 52.81, 84.965, 70.178, 69.185, 74.915, 82.202, 13.249, 
    82.25, 11.281, 93.171, 73.475, 90.46, 90.6, 0.52265, 87.431, 8.1774, 
    27.9, 42.096, 97.352, 79.064, 64.07, 2.1103, 8.4627, 68.265, 92.985, 
    50.946, 69.446, 7.1592, 24.182, 66.757, 57.598, 2.9508, 75.779, 0.047351, 
    41.469, 76.356, 61.54, 93.246, 25.649, 45.044, 24.801, 50.286, 79.97, 
    59.547, 93.619, 41.203, 21.246, 43.414, 0.45876, 42.524, 20.15, 84.761, 
    23.626, 48.619, 44.836, 82.783, 57.025, 41.581, 51.194, 71.778, 53.098, 
    72.192, 60.728, 15.655, 81.122, 19.691, 80.011, 57.605, 51.077, 80.47, 
    64.565 ;

 bangle_opt_qual =
  3.2595, 7.5256, 66.058, 88.903, 74.898, 76.374, 96.071, 13.906, 0.14014, 
    27.252, 18.001, 95.36, 57.473, 84.965, 83.568, 92.02, 13.609, 84.523, 
    58.668, 86.368, 45.412, 45.525, 8.6621, 30.995, 9.7682, 31.882, 81.59, 
    96.691, 65.721, 55.022, 1.1916, 18.689, 80.126, 9.2817, 0.85699, 23.315, 
    71.118, 34.074, 39.778, 12.915, 63.766, 64.981, 47.392, 59.783, 69.146, 
    55.591, 77.749, 59.256, 68.995, 47.61, 80.786, 58.156, 55.818, 14.701, 
    87.826, 17.311, 55.844, 52.687, 30.036, 85.658, 80.868, 52.541, 17.179, 
    85.649, 66.245, 75.881, 29.012, 41.347, 8.3909, 47.966, 35.914, 32.372, 
    39.492, 24.916, 34.734, 36.836, 19.52, 52.236, 43.165, 73.158, 65.935, 
    96.731, 71.646, 71.413, 78.351, 73.319, 46.687, 61.493, 85.207, 83.443, 
    2.4079, 46.688, 90.053, 18.48, 10.63, 62.944, 17.822, 52.88, 15.183, 
    67.028 ;

 alt_refrac =
  14587, 42597, 84486, 70892, 87112, 54446, 9280.7, 84977, 31139, 62813, 
    95070, 67686, 80786, 89199, 20464, 43174, 26857, 51477, 2412.6, 75411, 
    79259, 59639, 53438, 37797, 30940, 40733, 4017.5, 6242.5, 13729, 26045, 
    38100, 546.02, 53781, 46648, 51113, 72576, 76498, 75560, 9471.4, 21924, 
    31844, 80390, 89513, 25651, 87437, 40347, 1632, 43026, 65900, 80876, 
    89111, 22439, 50114, 74512, 50583, 76721, 29949, 94268, 90194, 78536, 
    92486, 73981, 48232, 35624, 53922, 3598, 11449, 64334, 94006, 12284, 
    51972, 5032, 60666, 58373, 88572, 84609, 68838, 78583, 55634, 1895, 
    1583.6, 57679, 11919, 25102, 31654, 66951, 57544, 36997, 66949, 29076, 
    88823, 53724, 41269, 84881, 41940, 42670, 69285, 85906, 62522, 42354 ;

 geop_refrac =
  37605, 78737, 63490, 27528, 10165, 53906, 5893.5, 40899, 56835, 71504, 
    68889, 93342, 30560, 68838, 46088, 22378, 44021, 16510, 50198, 97168, 
    49886, 91746, 53501, 70551, 43410, 24645, 75743, 6445.5, 5915.2, 61447, 
    97484, 39257, 53314, 61255, 65773, 57884, 24329, 3560.5, 46397, 33898, 
    23837, 35158, 56234, 77468, 74627, 13689, 46170, 62768, 27473, 34939, 
    16227, 38032, 19383, 86705, 29926, 91740, 7652.3, 32608, 61591, 86310, 
    14546, 51749, 44207, 11694, 48329, 76539, 97004, 22808, 86394, 6821.4, 
    80842, 34955, 30715, 22733, 35199, 70594, 89550, 27000, 12605, 68215, 
    59597, 13805, 38071, 49235, 74753, 50222, 11222, 65929, 53449, 35813, 
    83019, 18150, 85089, 64431, 87772, 77832, 24701, 73461, 1717.2, 26012 ;

 refrac =
  286.11, 109.56, 477.48, 180.5, 230.27, 29.038, 474.58, 465.79, 90.338, 
    146.25, 211.42, 397.89, 196.36, 312.61, 270.55, 113.6, 193.59, 363.57, 
    171.79, 130.77, 127.29, 135.95, 374.43, 317.64, 254.28, 395.32, 176.49, 
    85.083, 432.7, 296.74, 436.37, 450.95, 364.78, 208.38, 469.52, 387.3, 
    369.97, 174.62, 104.73, 107.24, 443.34, 351.49, 221.34, 362.12, 360.46, 
    171.66, 209.26, 335.35, 444.75, 30.122, 379.76, 53.696, 138.41, 320.98, 
    477.18, 239.2, 51.496, 440.76, 187.92, 1.6698, 69.199, 166.77, 137.5, 
    429.06, 321.1, 137.66, 106.47, 98.655, 350.66, 70.864, 129.49, 33.895, 
    434.95, 169.23, 275.09, 331.44, 50.771, 122.25, 197.8, 256.3, 34.814, 
    231.52, 462.48, 53.751, 477.28, 59.415, 287.39, 107.84, 290.19, 207.38, 
    477.72, 398.24, 487.96, 382.4, 318.16, 364.85, 202.13, 71.522, 208.98, 
    365.48 ;

 refrac_sigma =
  4.3775, 47.83, 0.89119, 7.8554, 9.1554, 34.39, 33.68, 12.698, 46.156, 
    44.633, 15.369, 7.7369, 7.8519, 5.2856, 48.159, 10.549, 20.425, 27.38, 
    39.204, 23.173, 23.876, 8.9563, 33.308, 34.734, 4.3527, 22.431, 42.669, 
    5.5453, 15.516, 42.607, 39.382, 26.313, 35.04, 27.023, 13.978, 20.444, 
    16.222, 26.843, 30.575, 8.5942, 11.406, 42.636, 40.417, 18.86, 43.317, 
    10.909, 19.12, 40.149, 1.2643, 27.178, 30.056, 21.316, 34.196, 39.556, 
    30.93, 44.027, 5.0548, 16.856, 7.4358, 43.107, 13.457, 43.765, 39.572, 
    8.1583, 41.776, 7.2361, 38.843, 3.0729, 19.701, 48.19, 23.929, 18.768, 
    0.064352, 9.7301, 30.856, 13.264, 34.584, 38.201, 38.155, 23.206, 37.073, 
    47.386, 2.2284, 0.29263, 17.364, 41.647, 33.36, 39.698, 8.5418, 44.851, 
    46.81, 14.069, 3.4355, 17.793, 31.613, 33.729, 26.838, 23.208, 2.1166, 
    45.011 ;

 refrac_qual =
  92.359, 19.369, 35.059, 74.102, 44.706, 25.131, 96.417, 50.546, 53.285, 
    32.692, 56.683, 62.727, 24.389, 50.359, 72.666, 32.736, 40.116, 68.608, 
    91.735, 52.518, 71.988, 65.71, 30.707, 7.6424, 48.348, 51.466, 9.8545, 
    10.035, 48.615, 32.672, 19.665, 0.66429, 15.904, 76.492, 8.403, 90.296, 
    46.583, 19.042, 60.101, 28.033, 16.708, 72.831, 56.977, 86.673, 1.2426, 
    67.908, 11.813, 23.065, 40.644, 22.545, 96.472, 77.41, 92.232, 77.074, 
    38.941, 6.2758, 20.611, 17.533, 86.039, 50.887, 24.327, 38.888, 13.663, 
    1.5075, 65.732, 41.432, 19.739, 49.626, 81.407, 65.639, 59.382, 24.974, 
    1.6183, 52.989, 66.92, 57.433, 0.34589, 41.018, 26.486, 72.086, 78.861, 
    81.34, 31.195, 89.432, 58.758, 11.465, 33.518, 11.306, 57.222, 24.712, 
    69.514, 26.216, 58.643, 32.155, 21.254, 11.502, 88.54, 46.914, 73.571, 
    72.664 ;

 dry_temp =
  212.18, 241.5, 307.97, 328.81, 218.97, 184.23, 223.71, 162.43, 271.66, 
    189.87, 253.21, 258.65, 232.98, 205.49, 179.91, 209.14, 199.54, 165.59, 
    324.7, 256.55, 329.71, 155.47, 316.32, 331.88, 309.76, 275.14, 293.46, 
    193.09, 195.19, 212.51, 240.78, 201.18, 220.64, 295.83, 304.44, 289.11, 
    280.47, 321.2, 189.9, 313.64, 206.68, 343.26, 165.76, 221.11, 250.44, 
    164.28, 307.91, 182.56, 248.8, 329.02, 221.7, 336.99, 326.49, 222.9, 
    345.76, 299.13, 175.34, 275.01, 160.14, 287.1, 287.93, 345.65, 342.87, 
    162.43, 199.15, 308.43, 230.3, 229.49, 259.93, 258.67, 255, 150.02, 
    193.05, 190.62, 177.46, 337.85, 294.25, 205.88, 216.95, 306.91, 284.05, 
    311.99, 213.82, 328.66, 214.98, 221.49, 325.49, 292, 249.07, 222.07, 
    203.23, 188.79, 342.7, 263.9, 208.28, 275.28, 340.99, 290.66, 263.1, 
    234.27 ;

 dry_temp_sigma =
  37.351, 0.47828, 19.453, 46.873, 34.167, 12.715, 25.371, 28.698, 19.733, 
    27.374, 48.438, 9.5867, 4.1336, 18.374, 21.584, 19.684, 30.94, 18.101, 
    29.205, 17.537, 35.94, 23.812, 32.431, 2.7338, 10.312, 17.945, 36.023, 
    47.562, 37.458, 8.93, 36.11, 16.651, 11.258, 8.7814, 31.374, 3.4903, 
    48.637, 36.348, 5.8166, 48.086, 27.124, 3.9544, 27.942, 2.7913, 33.241, 
    28.878, 43.664, 47.572, 24.206, 39.537, 9.628, 38.373, 47.609, 28.049, 
    40.876, 37.722, 47.393, 30.57, 30.619, 24.98, 46.652, 42.85, 31.843, 
    40.582, 7.1287, 23.231, 19.639, 36.743, 39.223, 47.408, 12.08, 43.896, 
    41.277, 22.432, 25.999, 28.736, 3.6713, 5.4817, 44.194, 17.261, 21.467, 
    17.851, 34.049, 22.413, 44.988, 32.317, 29.778, 40.153, 36.345, 22.442, 
    45.433, 15.504, 1.7025, 45.491, 44.847, 1.9794, 6.4634, 48.024, 27.201, 
    13.148 ;

 dry_temp_qual =
  34.105, 71.268, 91.856, 90.007, 10.471, 43.906, 41.38, 54.513, 34.416, 
    61.477, 38.8, 89.699, 92.128, 54.955, 91.591, 0.78182, 22.489, 68.834, 
    71.164, 82.264, 79.512, 61.729, 48.519, 18.965, 74.409, 32.489, 83.969, 
    3.9594, 19.609, 46.087, 42.835, 6.4133, 2.5496, 13.883, 0.50079, 16.751, 
    33.8, 25.165, 53.132, 24.63, 84.304, 18.942, 39.074, 44.19, 25.626, 
    76.738, 52.277, 85.92, 58.428, 47.76, 88.542, 9.3586, 66.25, 56.218, 
    1.7598, 1.8447, 29.236, 57.492, 16.083, 36.233, 12.004, 84.2, 94.816, 
    83.028, 29.782, 79.942, 63.406, 56.845, 62.258, 76.786, 84.055, 21.93, 
    60.845, 40.372, 1.2328, 82.207, 38.582, 28.315, 16.235, 30.902, 82.549, 
    13.66, 92.15, 92.322, 58.198, 17.444, 84.548, 19.607, 85.724, 88.376, 
    29.886, 26.892, 57.92, 24.641, 12.906, 35.877, 49.107, 57.953, 31.431, 
    29.993 ;

 geop =
  26365, 52234, 86519, 86296, 90274, 68428, 53320, 29554, 42269, 74295, 
    49550, 1865, 45455, 87168, 49797, 274.23, 9066.8, 73048, 55420, 79430, 
    41618, 12849, 43742, 11330, 60426, 57638, 56719, 9575.3, 49385, 65543, 
    36159, 67395, -323.01, 91470, 68902, 9389.5, 29931, 9498.4, 32124, 76887, 
    5046.3, 8757.2, 56158, 27649, 76584, 535.44, 29797, 80904, 38774, 55846, 
    82572, 44408, 43626, 50491, 83736, 83316, 33397, 22418, 93937, 75753, 
    27944, 70012, 15927, 82275, 93544, 28660, 26951, 17341, 13190, 55260, 
    6506.4, 52603, 66391, 68631, 62253, 74684, 80498, 69640, 80448, 91716, 
    5440, 23240, 46348, 3651.6, 37845, 51500, 45346, 2930.3, 69012, 11499, 
    42758, 80246, 87611, 7749.6, 90126, 83673, 24961, 70445, 67208, 69818 ;

 geop_sigma =
  134.15, 483.4, 144.88, 484.08, 107.79, 104.14, 485.37, 216.62, 127.8, 
    107.81, 369.06, 44.063, 104.45, 288.32, 337.29, 40.135, 195.23, 50.641, 
    53.658, 439.9, 465.48, 202.08, 210.49, 273.12, 268.64, 478.81, 107.44, 
    159.99, 146.77, 212.1, 434.7, 169.41, 465.95, 393.59, 64.18, 330.34, 
    428.32, 370.24, 420.83, 72.499, 245.44, 256.17, 437.66, 197.19, 439.48, 
    328.02, 463.33, 94.586, 280.6, 306.88, 5.0654, 385.05, 53.361, 12.331, 
    182.8, 218.69, 18.608, 164.6, 80.118, 451.25, 93.952, 269.63, 88.586, 
    34.947, 328.95, 430.23, 202.44, 368.46, 134.09, 156.37, 371.13, 138.23, 
    382.33, 252.7, 10.854, 439.05, 400.96, 343.15, 237.43, 239.47, 204.95, 
    210.87, 247.07, 434.68, 390.88, 351.34, 75.057, 385.23, 246.12, 253.32, 
    125.45, 355.74, 343.7, 343.51, 99.207, 272.4, 376.52, 487.71, 223.11, 
    369.09 ;

 press =
  986, 153.1, 761.84, 34.486, 64.12, 104.78, 729.08, 1036.1, 770.82, 876.33, 
    205.19, 85.762, 737.19, 395.46, 178.29, 772, 706.37, 231.71, 1021, 377.2, 
    802.21, 547.32, 305.84, 921.29, 412.79, 289.41, 257.04, 912.05, 606.48, 
    522.07, 513.8, 706.16, 126.17, 454.87, 456.25, 433.14, 147.78, 949.43, 
    492.81, 478.92, 867.56, 1055, 480.48, 372.28, 831.9, 836.77, 848.96, 
    201.55, 494.67, 574.5, 721.66, 178.38, 1035.5, 843.65, 115.84, 860.87, 
    628.69, 333.91, 490.88, 474.85, 1059.4, 624.71, 1060.9, 1074.4, 857.59, 
    774.91, 664.33, 882.68, 210.4, 974.78, 198.84, 836.64, 792.77, 1042.3, 
    478.47, 14.178, 189.37, 292.85, 592.73, 716.15, 1028, 807.11, 615.14, 
    655.41, 178.87, 928.05, 328.41, 663.01, 718.53, 881.2, 991.65, 478.15, 
    600.87, 115.01, 543.38, 773.31, 882.5, 774.96, 652.53, 413.85 ;

 press_sigma =
  1.2335, 0.88562, 4.211, 0.17029, 3.3604, 0.88735, 1.9804, 2.9192, 4.0274, 
    3.3961, 4.6171, 1.4506, 2.2938, 4.8035, 3.1024, 1.922, 4.214, 0.37175, 
    1.194, 3.0282, 0.87881, 1.261, 2.0133, 0.89182, 0.38758, 3.383, 2.4006, 
    3.8358, 3.8233, 0.53557, 1.9629, 0.95736, 2.7578, 3.4398, 1.0571, 1.1762, 
    2.6575, 2.3697, 1.6959, 2.1628, 2.429, 4.2952, 0.65071, 2.2782, 0.055026, 
    2.6149, 0.89839, 1.9349, 2.5771, 2.8629, 3.8683, 2.9382, 2.731, 4.2034, 
    4.8281, 3.067, 3.8704, 2.5649, 1.5088, 1.1948, 4.5475, 4.4132, 1.4843, 
    2.4535, 0.45878, 0.92111, 2.5262, 3.0932, 1.9342, 0.21118, 4.6962, 
    3.1714, 4.6039, 2.0873, 0.0068349, 1.2664, 4.3132, 2.1824, 1.1602, 
    1.5589, 4.7455, 0.63538, 0.96734, 4.1259, 4.1134, 0.95253, 0.24747, 
    1.6775, 3.2918, 1.2527, 2.5739, 3, 2.4956, 3.572, 4.0405, 0.92284, 
    1.9165, 3.5698, 2.4557, 4.1936 ;

 temp =
  330.48, 326.42, 320.1, 237.06, 279.92, 216.93, 278.82, 291.75, 209.02, 
    215.13, 195.09, 237.36, 341.86, 333.77, 232.63, 313.5, 247.48, 276.07, 
    335.73, 222.79, 243.96, 246.27, 205.34, 266.77, 258, 181.52, 198.82, 
    327.25, 202.27, 183.4, 270.04, 201.25, 254.03, 318.78, 194.12, 236.06, 
    243.08, 326.93, 340.09, 297.8, 224.18, 317.02, 245.89, 252.86, 190.58, 
    166.52, 238.5, 292.22, 243.61, 294.36, 270.59, 328.17, 310.55, 262.99, 
    225.77, 163.57, 173.43, 255.23, 296.65, 337.41, 331.3, 174.06, 153.81, 
    238.28, 207.7, 165.6, 314.67, 196.44, 264.56, 283.28, 174.87, 178.74, 
    177.49, 233.04, 328.88, 244.47, 225.87, 219.28, 180.83, 216.65, 189.81, 
    234.83, 160.85, 236.68, 244.86, 335.53, 198.19, 327.63, 174.36, 202.94, 
    314.37, 203.01, 217.26, 236.27, 293.14, 236.67, 292.82, 303.67, 287.96, 
    300.66 ;

 temp_sigma =
  3.434, 3.0203, 0.21276, 3.2949, 4.4136, 0.77893, 4.4517, 3.7608, 2.8213, 
    4.4699, 0.054439, 2.0844, 3.9621, 2.0606, 2.0744, 0.80266, 2.6031, 
    0.78364, 0.3023, 0.40433, 1.9054, 2.1229, 4.2816, 2.7783, 1.3566, 1.3565, 
    4.1325, 1.6448, 2.0428, 2.1845, 1.6158, 2.8438, 1.114, 3.9926, 2.0725, 
    2.386, 0.88583, 4.2568, 3.7298, 2.2886, 3.092, 0.36703, 3.0091, 2.8874, 
    3.5833, 1.6767, 1.162, 1.362, 3.2137, 3.4843, 1.6698, 1.2527, 4.4071, 
    0.55405, 4.6222, 4.7005, 0.10546, 0.59368, 0.20221, 1.9754, 0.98789, 
    2.9027, 0.33854, 4.6183, 1.5744, 4.6034, 3.5291, 1.5508, 2.1954, 1.4222, 
    0.47782, 0.98105, 2.6176, 4.3936, 3.6278, 0.75118, 1.1897, 0.84408, 
    2.3645, 0.99296, 3.3833, 3.3439, 3.7404, 0.6569, 3.8102, 0.26659, 3.6684, 
    3.6409, 1.8164, 1.2623, 0.04296, 0.61858, 1.5232, 3.7638, 3.1449, 2.07, 
    0.25998, 4.5317, 1.3469, 3.1905 ;

 shum =
  39.663, 32.77, 21.832, 7.2084, 3.5141, 28.842, 31.996, 40.08, 0.4779, 
    29.916, 34.782, 6.7626, 6.5878, 21.157, 19.244, 40.494, 15.695, 28.631, 
    34.717, 36.729, 31.716, 32.072, 41.267, 25.133, 30.593, 2.1429, 24.193, 
    20.811, 0.19864, 39.593, 2.3307, 44.878, 21.216, 21.162, 35.936, 11.856, 
    46.696, 21.717, 18.378, 42.435, 32.987, 3.1179, 44.798, 34.406, 35.651, 
    29.675, 1.6991, 17.55, 44.361, 19.445, 39.341, 34.85, 7.446, 39.642, 
    12.595, 8.2536, 12.04, 1.798, 2.067, 8.2414, 31.042, 45.244, 8.502, 
    34.557, 29.578, 2.5045, 31.246, 35.398, 11.065, 23.204, 28.567, 11.472, 
    38.04, 42.119, 33.578, 34.482, 45.991, 9.6555, 13.884, 6.3228, 30.5, 
    35.028, 5.046, 15.487, 43.9, 32.321, 3.0711, 38.879, 40.854, 5.3422, 
    2.8727, 19.891, 41.67, 29.903, 35.752, 23.873, 4.7724, 36.397, 13.714, 
    40.292 ;

 shum_sigma =
  2.879, 1.4039, 4.4724, 3.9166, 3.928, 4.3804, 0.57901, 3.2788, 0.20298, 
    4.5818, 2.7476, 4.668, 1.1956, 2.2539, 2.2449, 2.9525, 2.5029, 4.1193, 
    0.26739, 3.7394, 3.5276, 2.1644, 2.3975, 0.27867, 1.3924, 0.71069, 
    0.40326, 4.2303, 0.14769, 0.532, 2.1114, 1.4149, 2.9349, 1.3769, 0.85083, 
    4.1469, 3.2512, 0.98503, 4.8265, 2.2769, 0.92544, 2.6622, 2.9596, 3.9746, 
    3.2789, 4.0314, 1.563, 4.7205, 3.5068, 1.9441, 4.6258, 3.5596, 2.5869, 
    3.174, 2.1058, 3.0323, 3.0067, 0.55205, 1.0313, 1.3125, 1.9751, 4.0087, 
    0.90567, 0.25757, 1.4475, 3.4461, 1.1526, 3.3582, 4.2656, 4.4323, 1.2296, 
    2.2407, 3.6574, 1.3419, 0.65045, 1.0579, 2.4097, 0.28098, 2.5563, 2.8884, 
    1.382, 2.3292, 2.1914, 0.35576, 1.7965, 3.639, 1.4718, 4.012, 2.1559, 
    0.90484, 2.2166, 3.5365, 2.7951, 2.7957, 0.223, 2.1497, 4.1217, 3.9337, 
    4.8363, 3.4153 ;

 meteo_qual =
  28.79, 88.362, 26.604, 40.253, 25.138, 95.597, 24.255, 44.718, 86.398, 
    54.927, 58.625, 23.397, 66.785, 66.178, 27.501, 34.465, 11.839, 35.972, 
    95.299, 11.459, 77.356, 63.084, 55.441, 46.287, 12.949, 36.452, 19.499, 
    32.461, 6.239, 57.039, 51.412, 49.761, 74.22, 9.4576, 55.161, 76.774, 
    5.5672, 57.742, 16.338, 2.2382, 17.689, 10.165, 73.957, 67.596, 27.947, 
    45.408, 40.065, 90.025, 53.061, 26.9, 72.223, 29.363, 29.268, 94.373, 
    4.9978, 53.623, 56.474, 75.789, 86.417, 96.217, 94.15, 5.9706, 2.3335, 
    33.988, 60.851, 86.009, 82.361, 23.7, 59.543, 47.575, 3.6158, 14.217, 
    58.19, 64.003, 65.362, 25.252, 6.9485, 0.76631, 31.915, 36.688, 33.823, 
    47.266, 31.143, 51.756, 70.541, 28.933, 63.052, 92.507, 9.0377, 86.422, 
    89.927, 15.441, 93.51, 68.825, 50.837, 25.713, 16.831, 35.218, 33.981, 
    84.029 ;

 geop_sfc = 9549.3 ;

 press_sfc = 271.16 ;

 press_sfc_sigma = 1.6328 ;

 press_sfc_qual = 67.21 ;

 tph_bangle = 6.5714e+06 ;

 tpa_bangle = 0.0023606 ;

 tph_bangle_flag = 245 ;

 tph_refrac = 30056 ;

 tpn_refrac = 232.77 ;

 tph_refrac_flag = 179 ;

 tph_tdry_lrt = 27838 ;

 tpt_tdry_lrt = 279.23 ;

 tph_tdry_lrt_flag = 124 ;

 tph_tdry_cpt = 63756 ;

 tpt_tdry_cpt = 199.74 ;

 tph_tdry_cpt_flag = 240 ;

 prh_tdry_cpt = 90451 ;

 prt_tdry_cpt = 251.75 ;

 prh_tdry_cpt_flag = 44 ;

 tph_temp_lrt = 73654 ;

 tpt_temp_lrt = 220.14 ;

 tph_temp_lrt_flag = 89 ;

 tph_temp_cpt = 57660 ;

 tpt_temp_cpt = 292.63 ;

 tph_temp_cpt_flag = 31 ;

 prh_temp_cpt = 59330 ;

 prt_temp_cpt = 167.31 ;

 prh_temp_cpt_flag = 203 ;

 level_type =
  "HIRLAM" ;

 level_coeff_a =
  918.44, 478.52, 49.153, 1817.3, 346.28, 292.82, 1574.9, 1834.5, 1038.3, 
    52.552, 1383.2, 697.4, 1941.9, 1716, 1040.9, 542.62, 1939.3, 1258, 
    780.86, 1803.5, 356.99, 643.4, 1785.3, 389.08, 1754.2, 252.08, 773.3, 
    741.09, 981.82, 1097.2, 925.91, 1430.2, 421.54, 1688.3, 1079.2, 1112.8, 
    1880.8, 877.37, 963.91, 1860, 149.42, 1879.9, 867.78, 38.081, 1303.5, 
    332.05, 517.08, 1570.6, 792.12, 73.288, 381.11, 1755.9, 1885.1, 1856.4, 
    705.18, 1865.1, 1204.4, 1691, 365.41, 773.05, 1018.5, 1229, 1628.9, 
    1173.2, 889.96, 54.723, 294, 1222.3, 979.87, 493.67, 293.51, 1840.5, 
    272.09, 1392.6, 1376.3, 437.54, 1258.5, 1074.7, 836.13, 1711.4, 1580.9, 
    859.59, 664.55, 654.36, 933.32, 937.13, 823.15, 306.77, 434.2, 318.81, 
    1771.5, 564.94, 1382.1, 390.16, 1047.9, 760.62, 828.1, 1105.8, 801.95, 
    1190 ;

 level_coeff_b =
  0.60201, 1.858, 0.77243, 0.77784, 0.37778, 1.9429, 1.6231, 0.71016, 
    0.80909, 1.9235, 1.0144, 1.2078, 1.2836, 1.3377, 1.6191, 0.63902, 1.8711, 
    0.97076, 0.61386, 0.040326, 0.87269, 0.74514, 0.32178, 1.0901, 1.6028, 
    1.0478, 1.0169, 1.4188, 1.4157, 0.33166, 0.86977, 0.5844, 1.6287, 1.8809, 
    0.36231, 1.31, 0.77211, 0.38452, 0.073173, 1.4213, 0.43925, 0.054162, 
    1.3255, 0.077696, 1.7722, 0.20472, 1.3063, 0.50494, 0.39611, 0.44918, 
    0.82111, 0.77282, 0.37721, 0.37342, 0.98512, 1.028, 0.16771, 0.17447, 
    1.103, 0.95456, 1.1754, 1.1923, 1.3776, 0.97507, 1.5139, 1.7785, 1.5685, 
    1.8445, 0.52652, 1.494, 0.97305, 0.5427, 0.9659, 0.25601, 1.6377, 
    0.27167, 0.22897, 1.5983, 1.3589, 1.5987, 0.64753, 1.8779, 0.033427, 
    0.2982, 0.057199, 0.22915, 1.0707, 1.0473, 0.58905, 0.55516, 1.0915, 
    1.3443, 1.3672, 1.3209, 0.71486, 1.9329, 0.33015, 0.31614, 0.48086, 
    0.68984 ;
}
