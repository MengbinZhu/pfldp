netcdf ropp_test2d {
dimensions:
	dim_unlim = UNLIMITED ; // (1 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1b = 250 ;
	dim_lev2b = 91 ;
	dim_horiz = 31 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 359.9 ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 359.9 ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float geop(dim_unlim, dim_horiz, dim_lev2b) ;
		geop:long_name = "Geopotential height above geoid for P,T,H" ;
		geop:units = "geopotential metres" ;
		geop:valid_range = -1000., 1.e+05 ;
	float geop_sigma(dim_unlim, dim_horiz, dim_lev2b) ;
		geop_sigma:long_name = "Estimated error (1-sigma) for geopotential height" ;
		geop_sigma:units = "geopotential metres" ;
		geop_sigma:valid_range = 0., 500. ;
	double press(dim_unlim, dim_horiz, dim_lev2b) ;
		press:long_name = "Pressure" ;
		press:units = "hPa" ;
		press:valid_range = 0.01, 1100. ;
	float press_sigma(dim_unlim, dim_horiz, dim_lev2b) ;
		press_sigma:long_name = "Estimated error (1-sigma) for pressure" ;
		press_sigma:units = "hPa" ;
		press_sigma:valid_range = 0., 5. ;
	double temp(dim_unlim, dim_horiz, dim_lev2b) ;
		temp:long_name = "Temperature" ;
		temp:units = "kelvin" ;
		temp:valid_range = 150., 350. ;
	float temp_sigma(dim_unlim, dim_horiz, dim_lev2b) ;
		temp_sigma:long_name = "Estimated error (1-sigma) for temperature" ;
		temp_sigma:units = "kelvin" ;
		temp_sigma:valid_range = 0., 5. ;
	double shum(dim_unlim, dim_horiz, dim_lev2b) ;
		shum:long_name = "Specific humidity" ;
		shum:units = "gram / kilogram" ;
		shum:valid_range = 0., 50. ;
	float shum_sigma(dim_unlim, dim_horiz, dim_lev2b) ;
		shum_sigma:long_name = "Estimated  error (1-sigma) in specific humidity" ;
		shum_sigma:units = "gram / kilogram" ;
		shum_sigma:valid_range = 0., 5. ;
	float meteo_qual(dim_unlim, dim_horiz, dim_lev2b) ;
		meteo_qual:long_name = "Quality value for meteorological data" ;
		meteo_qual:units = "percent" ;
		meteo_qual:valid_range = 0., 100. ;

// global attributes:
		:title = "Atmospheric background data for ROPP Radio Occultation data" ;
		:institution = "NONE" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "UNKNOWN" ;
		:processing_date = "9999-99-99 99:99:99.999" ;
		:pod_method = "UNKNOWN" ;
		:phase_method = "UNKNOWN" ;
		:bangle_method = "UNKNOWN" ;
		:refrac_method = "UNKNOWN" ;
		:meteo_method = "UNKNOWN" ;
		:thin_method = "UNKNOWN" ;
		:software_version = "UNKNOWN" ;
data:

 occ_id =
  "OC_99999999999999_UNKN_U999_UNKN" ;

 gns_id =
  "U999" ;

 leo_id =
  "UNKN" ;

 stn_id =
  "UNKN" ;

 start_time = 0 ;

 year = 9999 ;

 month = 99 ;

 day = 99 ;

 hour = 99 ;

 minute = 99 ;

 second = 99 ;

 msec = 999 ;

 pcd = 65535 ;

 overall_qual = -9.9999e+07 ;

 time = 0 ;

 time_offset = 0 ;

 lat = -5.2 ;

 lon = -8.15 ;

 undulation = 10 ;

 roc = 6.371e+06 ;

 r_coc =
  0, 0, 0 ;

 azimuth = 1.05 ;

 lat_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 lon_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 azimuth_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 impact_L1 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 impact_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 impact =
  6.3737e+06, 6.3739e+06, 6.3741e+06, 6.3743e+06, 6.3745e+06, 6.3747e+06, 
    6.3749e+06, 6.3751e+06, 6.3753e+06, 6.3755e+06, 6.3757e+06, 6.3759e+06, 
    6.3761e+06, 6.3763e+06, 6.3765e+06, 6.3767e+06, 6.3769e+06, 6.3771e+06, 
    6.3773e+06, 6.3775e+06, 6.3777e+06, 6.3779e+06, 6.3781e+06, 6.3783e+06, 
    6.3785e+06, 6.3787e+06, 6.3789e+06, 6.3791e+06, 6.3793e+06, 6.3795e+06, 
    6.3797e+06, 6.3799e+06, 6.3801e+06, 6.3803e+06, 6.3805e+06, 6.3807e+06, 
    6.3809e+06, 6.3811e+06, 6.3813e+06, 6.3815e+06, 6.3817e+06, 6.3819e+06, 
    6.3821e+06, 6.3823e+06, 6.3825e+06, 6.3827e+06, 6.3829e+06, 6.3831e+06, 
    6.3833e+06, 6.3835e+06, 6.3837e+06, 6.3839e+06, 6.3841e+06, 6.3843e+06, 
    6.3845e+06, 6.3847e+06, 6.3849e+06, 6.3851e+06, 6.3853e+06, 6.3855e+06, 
    6.3857e+06, 6.3859e+06, 6.3861e+06, 6.3863e+06, 6.3865e+06, 6.3867e+06, 
    6.3869e+06, 6.3871e+06, 6.3873e+06, 6.3875e+06, 6.3877e+06, 6.3879e+06, 
    6.3881e+06, 6.3883e+06, 6.3885e+06, 6.3887e+06, 6.3889e+06, 6.3891e+06, 
    6.3893e+06, 6.3895e+06, 6.3897e+06, 6.3899e+06, 6.3901e+06, 6.3903e+06, 
    6.3905e+06, 6.3907e+06, 6.3909e+06, 6.3911e+06, 6.3913e+06, 6.3915e+06, 
    6.3917e+06, 6.3919e+06, 6.3921e+06, 6.3923e+06, 6.3925e+06, 6.3927e+06, 
    6.3929e+06, 6.3931e+06, 6.3933e+06, 6.3935e+06, 6.3937e+06, 6.3939e+06, 
    6.3941e+06, 6.3943e+06, 6.3945e+06, 6.3947e+06, 6.3949e+06, 6.3951e+06, 
    6.3953e+06, 6.3955e+06, 6.3957e+06, 6.3959e+06, 6.3961e+06, 6.3963e+06, 
    6.3965e+06, 6.3967e+06, 6.3969e+06, 6.3971e+06, 6.3973e+06, 6.3975e+06, 
    6.3977e+06, 6.3979e+06, 6.3981e+06, 6.3983e+06, 6.3985e+06, 6.3987e+06, 
    6.3989e+06, 6.3991e+06, 6.3993e+06, 6.3995e+06, 6.3997e+06, 6.3999e+06, 
    6.4001e+06, 6.4003e+06, 6.4005e+06, 6.4007e+06, 6.4009e+06, 6.4011e+06, 
    6.4013e+06, 6.4015e+06, 6.4017e+06, 6.4019e+06, 6.4021e+06, 6.4023e+06, 
    6.4025e+06, 6.4027e+06, 6.4029e+06, 6.4031e+06, 6.4033e+06, 6.4035e+06, 
    6.4037e+06, 6.4039e+06, 6.4041e+06, 6.4043e+06, 6.4045e+06, 6.4047e+06, 
    6.4049e+06, 6.4051e+06, 6.4053e+06, 6.4055e+06, 6.4057e+06, 6.4059e+06, 
    6.4061e+06, 6.4063e+06, 6.4065e+06, 6.4067e+06, 6.4069e+06, 6.4071e+06, 
    6.4073e+06, 6.4075e+06, 6.4077e+06, 6.4079e+06, 6.4081e+06, 6.4083e+06, 
    6.4085e+06, 6.4087e+06, 6.4089e+06, 6.4091e+06, 6.4093e+06, 6.4095e+06, 
    6.4097e+06, 6.4099e+06, 6.4101e+06, 6.4103e+06, 6.4105e+06, 6.4107e+06, 
    6.4109e+06, 6.4111e+06, 6.4113e+06, 6.4115e+06, 6.4117e+06, 6.4119e+06, 
    6.4121e+06, 6.4123e+06, 6.4125e+06, 6.4127e+06, 6.4129e+06, 6.4131e+06, 
    6.4133e+06, 6.4135e+06, 6.4137e+06, 6.4139e+06, 6.4141e+06, 6.4143e+06, 
    6.4145e+06, 6.4147e+06, 6.4149e+06, 6.4151e+06, 6.4153e+06, 6.4155e+06, 
    6.4157e+06, 6.4159e+06, 6.4161e+06, 6.4163e+06, 6.4165e+06, 6.4167e+06, 
    6.4169e+06, 6.4171e+06, 6.4173e+06, 6.4175e+06, 6.4177e+06, 6.4179e+06, 
    6.4181e+06, 6.4183e+06, 6.4185e+06, 6.4187e+06, 6.4189e+06, 6.4191e+06, 
    6.4193e+06, 6.4195e+06, 6.4197e+06, 6.4199e+06, 6.4201e+06, 6.4203e+06, 
    6.4205e+06, 6.4207e+06, 6.4209e+06, 6.4211e+06, 6.4213e+06, 6.4215e+06, 
    6.4217e+06, 6.4219e+06, 6.4221e+06, 6.4223e+06, 6.4225e+06, 6.4227e+06, 
    6.4229e+06, 6.4231e+06, 6.4233e+06, 6.4235e+06 ;

 impact_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 geop =
  10.389, 35.526, 70.442, 116.46, 173.6, 241.03, 320.25, 413.8, 522.3, 
    646.09, 785.65, 941.48, 1114, 1303.2, 1509.1, 1735.6, 1982.9, 2247.7, 
    2530.3, 2830.9, 3149.3, 3485.2, 3838.9, 4211.1, 4602.2, 5011.9, 5438.4, 
    5878.6, 6329.2, 6785.2, 7242.3, 7697.4, 8149.3, 8597.5, 9041.2, 9480.8, 
    9916.5, 10348, 10774, 11198, 11618, 12035, 12448, 12858, 13264, 13667, 
    14064, 14457, 14846, 15233, 15619, 16010, 16407, 16813, 17232, 17666, 
    18120, 18600, 19106, 19642, 20212, 20813, 21442, 22104, 22802, 23543, 
    24333, 25177, 26074, 27021, 28022, 29089, 30235, 31464, 32781, 34190, 
    35692, 37326, 39138, 41147, 43345, 45706, 48281, 51135, 54254, 57568, 
    61052, 64710, 68525, 72499, 78807,
  10.28, 35.414, 70.327, 116.34, 173.47, 240.9, 320.1, 413.64, 522.12, 645.9, 
    785.45, 941.26, 1113.8, 1302.9, 1508.9, 1735.4, 1982.7, 2247.4, 2529.9, 
    2830.5, 3148.8, 3484.7, 3838.4, 4210.7, 4601.9, 5011.7, 5438.1, 5878.5, 
    6329.2, 6785.2, 7242.2, 7697.2, 8149.1, 8597.1, 9040.8, 9480.4, 9916, 
    10347, 10774, 11197, 11617, 12034, 12447, 12857, 13263, 13666, 14063, 
    14456, 14845, 15232, 15619, 16009, 16406, 16813, 17231, 17666, 18120, 
    18599, 19105, 19641, 20211, 20812, 21442, 22104, 22803, 23542, 24332, 
    25177, 26074, 27021, 28021, 29088, 30235, 31462, 32778, 34188, 35692, 
    37328, 39137, 41144, 43343, 45706, 48281, 51135, 54254, 57569, 61052, 
    64709, 68524, 72500, 78809,
  10.268, 35.411, 70.335, 116.36, 173.52, 240.96, 320.2, 413.77, 522.29, 
    646.11, 785.69, 941.53, 1114, 1303.1, 1509.2, 1735.7, 1982.8, 2247.5, 
    2530, 2830.4, 3148.7, 3484.5, 3838.3, 4210.7, 4602, 5011.6, 5438, 5878.6, 
    6329.4, 6785.4, 7242.3, 7697.2, 8148.9, 8596.9, 9040.6, 9480.2, 9915.7, 
    10347, 10774, 11197, 11616, 12033, 12446, 12856, 13262, 13665, 14063, 
    14456, 14845, 15232, 15619, 16009, 16405, 16812, 17231, 17666, 18120, 
    18598, 19104, 19640, 20210, 20812, 21442, 22105, 22803, 23542, 24332, 
    25177, 26074, 27020, 28020, 29088, 30235, 31462, 32776, 34186, 35693, 
    37330, 39136, 41140, 43342, 45707, 48281, 51134, 54254, 57570, 61052, 
    64709, 68524, 72500, 78811,
  10.352, 35.506, 70.446, 116.49, 173.67, 241.15, 320.42, 414.04, 522.61, 
    646.48, 786.11, 941.99, 1114.5, 1303.6, 1509.7, 1736.2, 1983.3, 2247.8, 
    2530.3, 2830.6, 3148.8, 3484.6, 3838.4, 4210.9, 4602.1, 5011.6, 5438.2, 
    5879, 6329.9, 6785.8, 7242.7, 7697.5, 8149.2, 8597, 9040.7, 9480.3, 
    9915.8, 10347, 10774, 11197, 11616, 12032, 12446, 12855, 13262, 13664, 
    14062, 14456, 14846, 15233, 15619, 16008, 16405, 16811, 17231, 17666, 
    18120, 18597, 19103, 19639, 20210, 20812, 21443, 22105, 22804, 23543, 
    24332, 25177, 26074, 27020, 28019, 29087, 30235, 31461, 32775, 34185, 
    35694, 37333, 39136, 41137, 43340, 45708, 48282, 51134, 54254, 57571, 
    61053, 64709, 68524, 72499, 78811,
  10.41, 35.585, 70.556, 116.64, 173.88, 241.42, 320.77, 414.48, 523.17, 
    647.19, 786.99, 943.04, 1115.6, 1304.8, 1511.1, 1737.3, 1984, 2248.7, 
    2531.1, 2831.3, 3149.4, 3485.1, 3838.9, 4211.3, 4602.3, 5011.8, 5438.6, 
    5879.7, 6330.6, 6786.5, 7243.3, 7698.2, 8149.8, 8597.6, 9041.3, 9480.8, 
    9916.2, 10347, 10774, 11197, 11616, 12032, 12445, 12855, 13261, 13664, 
    14062, 14456, 14846, 15233, 15619, 16008, 16404, 16811, 17231, 17667, 
    18120, 18597, 19102, 19639, 20209, 20812, 21443, 22106, 22804, 23543, 
    24333, 25177, 26074, 27020, 28019, 29087, 30235, 31461, 32773, 34183, 
    35694, 37336, 39136, 41135, 43339, 45709, 48282, 51134, 54254, 57571, 
    61054, 64710, 68524, 72499, 78812,
  10.444, 35.645, 70.653, 116.79, 174.08, 241.7, 321.14, 414.96, 523.79, 
    647.97, 787.95, 944.15, 1116.8, 1306, 1512.3, 1738.3, 1984.8, 2249.4, 
    2531.8, 2832, 3149.9, 3485.6, 3839.4, 4211.7, 4602.5, 5012, 5439, 5880.3, 
    6331.2, 6787.1, 7244, 7698.8, 8150.4, 8598.2, 9041.8, 9481.1, 9916.4, 
    10347, 10774, 11197, 11616, 12032, 12445, 12855, 13261, 13663, 14062, 
    14456, 14846, 15233, 15619, 16008, 16403, 16810, 17231, 17667, 18120, 
    18596, 19102, 19638, 20209, 20812, 21443, 22107, 22805, 23543, 24333, 
    25178, 26074, 27019, 28018, 29087, 30235, 31461, 32772, 34181, 35695, 
    37339, 39137, 41133, 43338, 45710, 48283, 51133, 54253, 57571, 61055, 
    64711, 68525, 72499, 78812,
  10.469, 35.663, 70.662, 116.78, 174.06, 241.65, 321.06, 414.84, 523.62, 
    647.74, 787.68, 943.95, 1116.8, 1306.3, 1512.8, 1738.4, 1984.5, 2249.3, 
    2531.6, 2831.8, 3149.8, 3485.5, 3839.3, 4211.4, 4602.3, 5011.8, 5438.8, 
    5880.1, 6331, 6786.8, 7243.7, 7698.6, 8150.2, 8597.9, 9041.4, 9480.7, 
    9915.9, 10347, 10773, 11196, 11615, 12031, 12444, 12854, 13260, 13662, 
    14061, 14456, 14846, 15233, 15619, 16007, 16402, 16809, 17230, 17666, 
    18119, 18595, 19101, 19637, 20208, 20812, 21443, 22106, 22804, 23543, 
    24332, 25177, 26073, 27018, 28018, 29086, 30235, 31460, 32771, 34180, 
    35694, 37340, 39138, 41132, 43336, 45709, 48283, 51132, 54251, 57570, 
    61056, 64712, 68525, 72497, 78810,
  10.459, 35.644, 70.631, 116.74, 173.99, 241.56, 320.93, 414.67, 523.39, 
    647.45, 787.34, 943.67, 1116.7, 1306.5, 1513.3, 1738.4, 1984.1, 2249, 
    2531.3, 2831.6, 3149.6, 3485.4, 3839.1, 4211.3, 4602.1, 5011.7, 5438.8, 
    5880, 6330.8, 6786.5, 7243.3, 7698.2, 8149.8, 8597.5, 9041, 9480.2, 
    9915.3, 10346, 10773, 11195, 11614, 12030, 12443, 12853, 13259, 13661, 
    14060, 14455, 14845, 15233, 15619, 16007, 16401, 16807, 17229, 17665, 
    18118, 18594, 19100, 19637, 20208, 20811, 21443, 22106, 22804, 23542, 
    24332, 25177, 26072, 27017, 28017, 29086, 30234, 31458, 32770, 34178, 
    35694, 37341, 39138, 41131, 43333, 45708, 48283, 51131, 54249, 57570, 
    61057, 64713, 68525, 72495, 78809,
  10.45, 35.636, 70.622, 116.73, 173.98, 241.54, 320.91, 414.63, 523.34, 
    647.38, 787.26, 943.64, 1116.8, 1306.8, 1513.9, 1738.8, 1984.2, 2249.1, 
    2531.5, 2831.8, 3149.9, 3485.8, 3839.6, 4211.8, 4602.8, 5012.5, 5439.6, 
    5880.7, 6331.3, 6786.9, 7243.7, 7698.7, 8150.3, 8598, 9041.4, 9480.5, 
    9915.7, 10347, 10773, 11196, 11615, 12031, 12444, 12853, 13259, 13661, 
    14060, 14455, 14846, 15234, 15620, 16008, 16401, 16807, 17228, 17664, 
    18117, 18594, 19100, 19638, 20209, 20813, 21445, 22107, 22804, 23543, 
    24332, 25178, 26073, 27016, 28017, 29087, 30234, 31458, 32769, 34177, 
    35695, 37342, 39140, 41132, 43332, 45707, 48283, 51131, 54248, 57570, 
    61059, 64716, 68525, 72494, 78807,
  10.373, 35.564, 70.555, 116.67, 173.93, 241.5, 320.87, 414.61, 523.32, 
    647.37, 787.27, 943.71, 1117, 1307.2, 1514.5, 1739.3, 1984.4, 2249.3, 
    2531.7, 2832.1, 3150.4, 3486.4, 3840.1, 4212.4, 4603.5, 5013.3, 5440.5, 
    5881.5, 6331.8, 6787.3, 7244.1, 7699.2, 8150.8, 8598.4, 9041.8, 9480.9, 
    9916.1, 10347, 10774, 11196, 11615, 12031, 12444, 12853, 13259, 13661, 
    14060, 14455, 14846, 15234, 15621, 16009, 16401, 16806, 17228, 17664, 
    18117, 18593, 19100, 19638, 20210, 20814, 21446, 22108, 22804, 23543, 
    24333, 25178, 26073, 27016, 28018, 29088, 30234, 31457, 32769, 34177, 
    35695, 37343, 39141, 41133, 43331, 45707, 48284, 51131, 54248, 57571, 
    61062, 64718, 68526, 72492, 78806,
  10.296, 35.496, 70.5, 116.63, 173.91, 241.51, 320.92, 414.7, 523.47, 
    647.57, 787.55, 944.05, 1117.3, 1307.6, 1515, 1739.7, 1984.5, 2249.3, 
    2531.9, 2832.4, 3150.6, 3486.5, 3840.3, 4212.7, 4603.9, 5013.7, 5440.8, 
    5881.6, 6331.7, 6787.1, 7244, 7699.1, 8150.7, 8598.2, 9041.5, 9480.6, 
    9915.9, 10347, 10774, 11196, 11614, 12030, 12443, 12852, 13258, 13660, 
    14059, 14455, 14846, 15234, 15621, 16009, 16401, 16805, 17226, 17662, 
    18115, 18592, 19099, 19638, 20210, 20814, 21446, 22108, 22803, 23542, 
    24333, 25178, 26072, 27015, 28018, 29089, 30234, 31456, 32767, 34176, 
    35696, 37343, 39141, 41133, 43328, 45705, 48283, 51130, 54246, 57571, 
    61063, 64719, 68525, 72489, 78804,
  10.252, 35.459, 70.475, 116.62, 173.93, 241.56, 321, 414.82, 523.62, 
    647.79, 787.83, 944.37, 1117.7, 1308, 1515.4, 1740.1, 1984.7, 2249.4, 
    2532, 2832.6, 3150.9, 3486.7, 3840.4, 4212.8, 4604.2, 5014, 5441.1, 
    5881.7, 6331.5, 6786.9, 7244, 7699.1, 8150.6, 8597.9, 9041.1, 9480.2, 
    9915.6, 10347, 10773, 11195, 11614, 12030, 12443, 12852, 13257, 13659, 
    14059, 14454, 14846, 15234, 15622, 16009, 16401, 16804, 17224, 17660, 
    18113, 18590, 19098, 19639, 20211, 20814, 21447, 22108, 22802, 23541, 
    24332, 25178, 26072, 27014, 28017, 29089, 30233, 31454, 32765, 34175, 
    35696, 37343, 39141, 41132, 43325, 45702, 48282, 51128, 54245, 57571, 
    61065, 64720, 68524, 72486, 78802,
  10.322, 35.529, 70.547, 116.7, 174, 241.63, 321.07, 414.89, 523.7, 647.86, 
    787.91, 944.46, 1117.8, 1308.2, 1515.6, 1740.4, 1985.1, 2249.7, 2532.3, 
    2833, 3151.3, 3487.1, 3840.7, 4213.2, 4604.6, 5014.5, 5441.5, 5881.9, 
    6331.5, 6787, 7244.2, 7699.3, 8150.7, 8598, 9041, 9480.3, 9915.7, 10347, 
    10773, 11195, 11614, 12029, 12442, 12851, 13257, 13659, 14058, 14454, 
    14846, 15235, 15622, 16010, 16401, 16803, 17223, 17659, 18112, 18589, 
    19098, 19639, 20212, 20815, 21447, 22108, 22802, 23540, 24332, 25178, 
    26072, 27014, 28017, 29090, 30234, 31454, 32763, 34174, 35697, 37343, 
    39141, 41131, 43322, 45700, 48281, 51127, 54245, 57572, 61066, 64721, 
    68522, 72483, 78801,
  10.427, 35.627, 70.635, 116.77, 174.06, 241.66, 321.08, 414.86, 523.64, 
    647.76, 787.78, 944.31, 1117.7, 1308.1, 1515.6, 1740.6, 1985.3, 2249.9, 
    2532.5, 2833.2, 3151.6, 3487.4, 3841, 4213.3, 4604.8, 5014.8, 5441.6, 
    5881.9, 6331.4, 6786.9, 7244.3, 7699.4, 8150.7, 8597.8, 9040.8, 9480.1, 
    9915.6, 10347, 10773, 11195, 11613, 12029, 12442, 12851, 13256, 13658, 
    14058, 14454, 14846, 15235, 15623, 16010, 16401, 16802, 17221, 17657, 
    18110, 18588, 19097, 19640, 20212, 20815, 21447, 22107, 22801, 23540, 
    24332, 25178, 26071, 27013, 28017, 29091, 30234, 31453, 32762, 34173, 
    35697, 37343, 39141, 41131, 43319, 45697, 48280, 51126, 54244, 57573, 
    61068, 64721, 68520, 72480, 78800,
  10.441, 35.636, 70.634, 116.76, 174.03, 241.61, 321.01, 414.77, 523.51, 
    647.61, 787.65, 944.2, 1117.6, 1308.1, 1515.8, 1740.8, 1985.6, 2250.3, 
    2532.8, 2833.5, 3151.9, 3487.7, 3841.2, 4213.6, 4605.2, 5015.1, 5441.8, 
    5881.8, 6331.2, 6786.9, 7244.4, 7699.5, 8150.7, 8597.7, 9040.7, 9480.1, 
    9915.6, 10347, 10773, 11195, 11613, 12029, 12442, 12851, 13256, 13658, 
    14057, 14454, 14846, 15236, 15624, 16011, 16401, 16801, 17221, 17656, 
    18109, 18587, 19097, 19640, 20213, 20815, 21447, 22107, 22801, 23540, 
    24332, 25177, 26071, 27013, 28017, 29091, 30235, 31453, 32760, 34171, 
    35697, 37344, 39141, 41130, 43317, 45695, 48279, 51125, 54245, 57575, 
    61069, 64721, 68518, 72478, 78799,
  10.425, 35.616, 70.609, 116.73, 173.99, 241.57, 320.96, 414.71, 523.44, 
    647.55, 787.63, 944.23, 1117.7, 1308.3, 1516.1, 1741.2, 1986.1, 2250.7, 
    2533.3, 2834, 3152.4, 3488.2, 3841.6, 4214, 4605.8, 5015.8, 5442.2, 
    5881.9, 6331.2, 6787.1, 7244.8, 7699.8, 8150.9, 8597.8, 9040.8, 9480.3, 
    9915.8, 10347, 10773, 11195, 11613, 12029, 12442, 12851, 13256, 13658, 
    14058, 14454, 14847, 15237, 15625, 16012, 16401, 16801, 17220, 17656, 
    18109, 18587, 19097, 19640, 20213, 20815, 21447, 22107, 22801, 23540, 
    24333, 25177, 26070, 27013, 28017, 29092, 30236, 31453, 32759, 34171, 
    35697, 37344, 39142, 41131, 43315, 45692, 48277, 51124, 54246, 57576, 
    61070, 64721, 68516, 72476, 78799,
  10.396, 35.579, 70.562, 116.67, 173.92, 241.48, 320.85, 414.58, 523.28, 
    647.39, 787.5, 944.15, 1117.7, 1308.5, 1516.4, 1741.6, 1986.4, 2250.9, 
    2533.6, 2834.4, 3152.8, 3488.6, 3842.1, 4214.7, 4606.5, 5016.5, 5442.6, 
    5882, 6331.3, 6787.4, 7245.2, 7700.2, 8151.1, 8598, 9041.1, 9480.6, 
    9916.2, 10347, 10773, 11195, 11614, 12030, 12442, 12851, 13256, 13659, 
    14058, 14455, 14848, 15238, 15626, 16013, 16402, 16801, 17220, 17656, 
    18109, 18587, 19097, 19641, 20214, 20815, 21446, 22107, 22802, 23541, 
    24333, 25177, 26070, 27012, 28017, 29093, 30238, 31454, 32758, 34170, 
    35697, 37344, 39142, 41131, 43314, 45690, 48276, 51124, 54248, 57578, 
    61071, 64720, 68514, 72474, 78799,
  10.41, 35.575, 70.532, 116.6, 173.81, 241.31, 320.62, 414.29, 522.95, 
    647.05, 787.15, 943.85, 1117.5, 1308.3, 1516.3, 1741.7, 1986.3, 2250.6, 
    2533.3, 2834.1, 3152.7, 3488.6, 3842.2, 4214.9, 4606.8, 5016.6, 5442.3, 
    5881.4, 6330.6, 6787, 7244.9, 7699.7, 8150.6, 8597.4, 9040.7, 9480.3, 
    9915.7, 10346, 10773, 11195, 11613, 12029, 12442, 12851, 13256, 13658, 
    14058, 14454, 14848, 15238, 15626, 16014, 16402, 16801, 17219, 17655, 
    18108, 18586, 19096, 19640, 20214, 20815, 21445, 22106, 22801, 23541, 
    24333, 25176, 26068, 27011, 28016, 29093, 30238, 31454, 32756, 34169, 
    35696, 37343, 39142, 41131, 43312, 45686, 48273, 51123, 54250, 57580, 
    61070, 64717, 68510, 72471, 78798,
  10.451, 35.597, 70.528, 116.56, 173.72, 241.18, 320.43, 414.03, 522.64, 
    646.74, 786.85, 943.6, 1117.4, 1308.2, 1516.3, 1741.8, 1986.2, 2250.3, 
    2532.9, 2833.8, 3152.4, 3488.5, 3842.3, 4215, 4606.9, 5016.5, 5442, 
    5880.7, 6330.1, 6786.5, 7244.4, 7699.2, 8150, 8596.9, 9040.2, 9479.9, 
    9915.2, 10346, 10772, 11194, 11613, 12029, 12442, 12850, 13255, 13658, 
    14057, 14454, 14848, 15238, 15626, 16013, 16401, 16800, 17218, 17654, 
    18108, 18585, 19096, 19640, 20213, 20814, 21444, 22105, 22801, 23541, 
    24333, 25175, 26067, 27011, 28016, 29093, 30239, 31454, 32755, 34167, 
    35695, 37341, 39142, 41132, 43311, 45683, 48270, 51124, 54252, 57580, 
    61069, 64714, 68508, 72469, 78798,
  10.492, 35.622, 70.53, 116.54, 173.66, 241.08, 320.29, 413.84, 522.45, 
    646.56, 786.7, 943.53, 1117.4, 1308.3, 1516.5, 1742.1, 1986.4, 2250.1, 
    2532.7, 2833.6, 3152.3, 3488.5, 3842.5, 4215.3, 4607.1, 5016.7, 5442, 
    5880.6, 6330.1, 6786.7, 7244.6, 7699.3, 8150, 8597, 9040.5, 9480.2, 
    9915.5, 10346, 10772, 11195, 11614, 12030, 12442, 12850, 13255, 13658, 
    14058, 14455, 14848, 15239, 15627, 16014, 16402, 16800, 17218, 17654, 
    18108, 18586, 19096, 19640, 20214, 20814, 21444, 22105, 22801, 23542, 
    24333, 25175, 26067, 27011, 28017, 29094, 30240, 31454, 32755, 34167, 
    35694, 37340, 39142, 41134, 43311, 45680, 48268, 51126, 54255, 57582, 
    61068, 64712, 68506, 72468, 78798,
  10.528, 35.643, 70.531, 116.51, 173.61, 240.99, 320.16, 413.67, 522.27, 
    646.4, 786.58, 943.49, 1117.4, 1308.5, 1516.8, 1742.6, 1986.7, 2250, 
    2532.5, 2833.5, 3152.4, 3488.8, 3842.9, 4215.7, 4607.6, 5017.1, 5442.3, 
    5880.9, 6330.4, 6787.2, 7245.1, 7699.7, 8150.4, 8597.4, 9041.1, 9480.8, 
    9916.1, 10347, 10773, 11196, 11615, 12031, 12443, 12851, 13256, 13658, 
    14059, 14456, 14850, 15240, 15628, 16015, 16402, 16800, 17217, 17654, 
    18108, 18586, 19096, 19641, 20215, 20815, 21445, 22106, 22802, 23543, 
    24334, 25176, 26067, 27011, 28018, 29095, 30241, 31455, 32756, 34167, 
    35693, 37339, 39143, 41135, 43311, 45678, 48268, 51130, 54258, 57583, 
    61066, 64710, 68504, 72467, 78798,
  10.474, 35.595, 70.491, 116.48, 173.59, 241, 320.19, 413.73, 522.35, 
    646.47, 786.64, 943.52, 1117.4, 1308.5, 1516.8, 1742.7, 1986.7, 2249.7, 
    2532, 2833, 3152, 3488.4, 3842.6, 4215.5, 4607.3, 5016.8, 5441.9, 5880.6, 
    6330.3, 6787.1, 7244.9, 7699.4, 8150.1, 8597.2, 9040.9, 9480.6, 9915.8, 
    10347, 10773, 11196, 11615, 12031, 12443, 12851, 13255, 13658, 14058, 
    14456, 14849, 15240, 15628, 16014, 16402, 16799, 17216, 17653, 18107, 
    18586, 19096, 19640, 20214, 20815, 21444, 22105, 22802, 23543, 24334, 
    25175, 26066, 27011, 28018, 29094, 30240, 31455, 32756, 34167, 35691, 
    37337, 39143, 41136, 43310, 45675, 48268, 51133, 54260, 57582, 61063, 
    64707, 68502, 72466, 78797,
  10.38, 35.497, 70.388, 116.37, 173.48, 240.87, 320.05, 413.6, 522.21, 
    646.32, 786.47, 943.33, 1117.3, 1308.4, 1516.8, 1742.8, 1986.7, 2249.3, 
    2531.4, 2832.3, 3151.3, 3487.8, 3842, 4214.9, 4606.8, 5016.3, 5441.4, 
    5880.2, 6330.1, 6787, 7244.6, 7699, 8149.6, 8596.7, 9040.4, 9480, 9915.3, 
    10346, 10773, 11195, 11615, 12031, 12443, 12851, 13255, 13657, 14057, 
    14455, 14849, 15240, 15627, 16013, 16400, 16797, 17214, 17651, 18106, 
    18585, 19095, 19639, 20214, 20814, 21444, 22104, 22801, 23542, 24333, 
    25174, 26066, 27011, 28018, 29094, 30239, 31454, 32756, 34166, 35690, 
    37335, 39143, 41137, 43309, 45673, 48268, 51136, 54261, 57580, 61060, 
    64704, 68500, 72465, 78796,
  10.387, 35.497, 70.38, 116.35, 173.44, 240.82, 319.98, 413.49, 522.06, 
    646.11, 786.24, 943.09, 1117, 1308.2, 1516.7, 1742.8, 1986.8, 2249.2, 
    2530.9, 2831.7, 3150.7, 3487.3, 3841.6, 4214.6, 4606.6, 5016, 5441.1, 
    5880.1, 6330.3, 6787.2, 7244.8, 7699.1, 8149.6, 8596.8, 9040.5, 9480.1, 
    9915.4, 10346, 10773, 11196, 11615, 12031, 12443, 12851, 13255, 13657, 
    14057, 14455, 14849, 15240, 15628, 16014, 16400, 16797, 17214, 17651, 
    18106, 18584, 19095, 19639, 20214, 20815, 21444, 22105, 22801, 23543, 
    24333, 25174, 26066, 27011, 28018, 29094, 30238, 31454, 32757, 34167, 
    35689, 37334, 39144, 41138, 43309, 45672, 48271, 51140, 54262, 57579, 
    61057, 64702, 68499, 72465, 78796,
  10.501, 35.604, 70.477, 116.44, 173.51, 240.87, 320, 413.48, 521.99, 
    645.98, 786.09, 942.94, 1116.9, 1308.1, 1516.7, 1743, 1987, 2249.2, 
    2530.6, 2831.3, 3150.3, 3487, 3841.4, 4214.5, 4606.5, 5015.9, 5441.1, 
    5880.3, 6330.7, 6787.7, 7245.3, 7699.5, 8150, 8597.1, 9040.8, 9480.5, 
    9915.8, 10347, 10774, 11197, 11616, 12032, 12444, 12852, 13256, 13657, 
    14058, 14456, 14850, 15241, 15628, 16014, 16400, 16796, 17213, 17650, 
    18106, 18585, 19095, 19640, 20215, 20816, 21446, 22106, 22802, 23543, 
    24334, 25175, 26067, 27012, 28020, 29094, 30238, 31455, 32758, 34168, 
    35689, 37334, 39144, 41138, 43309, 45673, 48275, 51145, 54263, 57577, 
    61055, 64700, 68499, 72465, 78796,
  10.478, 35.585, 70.463, 116.43, 173.52, 240.88, 320.03, 413.52, 522.04, 
    646.04, 786.17, 943.03, 1117, 1308.2, 1516.8, 1743, 1987.1, 2249.4, 
    2530.6, 2831.2, 3150.1, 3486.7, 3841.1, 4214.3, 4606.1, 5015.5, 5440.9, 
    5880.2, 6330.8, 6787.9, 7245.4, 7699.6, 8150, 8597.2, 9040.9, 9480.5, 
    9915.8, 10347, 10774, 11197, 11616, 12033, 12445, 12852, 13256, 13657, 
    14057, 14455, 14850, 15241, 15628, 16014, 16400, 16796, 17212, 17649, 
    18105, 18584, 19095, 19639, 20215, 20817, 21446, 22106, 22802, 23543, 
    24333, 25175, 26067, 27013, 28020, 29095, 30237, 31454, 32758, 34168, 
    35689, 37333, 39144, 41138, 43310, 45674, 48278, 51147, 54262, 57575, 
    61053, 64700, 68499, 72464, 78796,
  10.412, 35.524, 70.409, 116.39, 173.48, 240.86, 320.02, 413.55, 522.08, 
    646.09, 786.23, 943.09, 1117.1, 1308.3, 1516.8, 1743, 1987.1, 2249.4, 
    2530.6, 2831, 3149.8, 3486.3, 3840.8, 4213.9, 4605.7, 5015.1, 5440.5, 
    5879.9, 6330.7, 6787.9, 7245.3, 7699.4, 8149.8, 8597, 9040.6, 9480.2, 
    9915.5, 10347, 10774, 11197, 11617, 12033, 12445, 12852, 13255, 13657, 
    14057, 14455, 14850, 15241, 15628, 16014, 16399, 16795, 17211, 17648, 
    18105, 18584, 19094, 19638, 20214, 20817, 21447, 22107, 22803, 23543, 
    24332, 25174, 26067, 27013, 28021, 29095, 30236, 31453, 32758, 34168, 
    35688, 37333, 39144, 41137, 43310, 45676, 48281, 51148, 54260, 57573, 
    61051, 64699, 68498, 72464, 78796,
  10.433, 35.547, 70.436, 116.42, 173.52, 240.91, 320.09, 413.64, 522.24, 
    646.29, 786.45, 943.31, 1117.3, 1308.5, 1517, 1743.2, 1987.2, 2249.5, 
    2530.8, 2831.1, 3149.8, 3486.3, 3840.8, 4214, 4605.7, 5015, 5440.4, 
    5879.9, 6330.7, 6787.9, 7245.3, 7699.3, 8149.8, 8596.9, 9040.6, 9480.1, 
    9915.4, 10347, 10774, 11197, 11617, 12033, 12445, 12852, 13255, 13656, 
    14056, 14454, 14849, 15241, 15628, 16014, 16399, 16794, 17210, 17648, 
    18104, 18584, 19094, 19638, 20214, 20817, 21448, 22107, 22803, 23542, 
    24332, 25174, 26067, 27013, 28021, 29096, 30236, 31452, 32759, 34169, 
    35689, 37333, 39143, 41135, 43310, 45678, 48283, 51149, 54259, 57571, 
    61050, 64698, 68499, 72464, 78796,
  10.485, 35.602, 70.495, 116.48, 173.59, 240.99, 320.17, 413.77, 522.43, 
    646.55, 786.73, 943.62, 1117.6, 1308.8, 1517.3, 1743.5, 1987.5, 2249.8, 
    2531.2, 2831.5, 3150.2, 3486.8, 3841.3, 4214.5, 4606.2, 5015.5, 5440.9, 
    5880.3, 6331.1, 6788.2, 7245.5, 7699.4, 8149.9, 8597.2, 9040.8, 9480.4, 
    9915.7, 10347, 10774, 11198, 11618, 12034, 12445, 12852, 13255, 13656, 
    14056, 14454, 14849, 15241, 15629, 16014, 16399, 16794, 17210, 17648, 
    18105, 18585, 19094, 19638, 20214, 20818, 21449, 22108, 22803, 23542, 
    24331, 25174, 26068, 27014, 28023, 29097, 30235, 31451, 32759, 34170, 
    35689, 37335, 39143, 41134, 43311, 45682, 48286, 51149, 54257, 57570, 
    61050, 64699, 68499, 72465, 78797,
  10.473, 35.598, 70.504, 116.51, 173.63, 241.05, 320.26, 413.87, 522.57, 
    646.73, 786.91, 943.8, 1117.8, 1308.9, 1517.4, 1743.6, 1987.6, 2250.1, 
    2531.5, 2831.8, 3150.5, 3487.2, 3841.8, 4215, 4606.7, 5016, 5441.4, 
    5880.7, 6331.4, 6788.3, 7245.5, 7699.3, 8149.9, 8597.2, 9040.9, 9480.4, 
    9915.8, 10347, 10774, 11198, 11618, 12034, 12446, 12853, 13256, 13656, 
    14055, 14454, 14849, 15241, 15629, 16014, 16399, 16794, 17210, 17648, 
    18105, 18585, 19094, 19638, 20215, 20819, 21449, 22109, 22803, 23541, 
    24331, 25174, 26068, 27015, 28024, 29097, 30235, 31451, 32759, 34170, 
    35690, 37336, 39143, 41132, 43312, 45685, 48287, 51147, 54256, 57569, 
    61050, 64699, 68500, 72465, 78798,
  10.497, 35.631, 70.545, 116.56, 173.7, 241.13, 320.36, 413.98, 522.68, 
    646.84, 787.01, 943.86, 1117.8, 1308.9, 1517.4, 1743.6, 1987.6, 2250.1, 
    2531.6, 2831.9, 3150.6, 3487.4, 3842.1, 4215.3, 4606.9, 5016.2, 5441.5, 
    5880.8, 6331.2, 6788, 7245, 7698.8, 8149.4, 8596.7, 9040.4, 9479.9, 
    9915.3, 10347, 10774, 11198, 11618, 12034, 12446, 12853, 13255, 13655, 
    14054, 14452, 14848, 15240, 15628, 16013, 16399, 16794, 17209, 17648, 
    18105, 18585, 19094, 19637, 20214, 20819, 21450, 22109, 22802, 23540, 
    24330, 25174, 26069, 27016, 28025, 29097, 30234, 31450, 32759, 34169, 
    35689, 37338, 39143, 41129, 43312, 45688, 48287, 51145, 54255, 57568, 
    61050, 64700, 68500, 72465, 78798 ;

 geop_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 press =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 947.06, 779.88, 634.17, 508.6, 
    401.76, 312.09, 238, 177.81, 129.85, 92.442, 63.957, 42.85, 27.683, 
    17.161, 10.148, 5.684, 2.9904, 1.015 ;

 press_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 temp =
  297.08, 296.78, 296.42, 295.96, 295.39, 294.73, 293.96, 293.05, 292, 290.8, 
    289.46, 288, 287, 285.14, 283.76, 291.72, 289.28, 287.36, 285.8, 283.73, 
    281.45, 279.32, 277.48, 276.07, 274.69, 272.98, 270.77, 268.83, 266.35, 
    263.35, 260.66, 257.36, 253.98, 250.14, 246.2, 242.7, 238.97, 235.04, 
    231.43, 228.52, 225.66, 222.46, 219.24, 216.05, 212.89, 209.43, 205.63, 
    202.07, 199.48, 197.59, 196.6, 196.94, 197.43, 197.5, 198.49, 199.76, 
    201.87, 204.4, 205.2, 208.69, 211.95, 211.5, 211.74, 212.5, 213.63, 
    216.38, 219.73, 222.46, 223.34, 222.62, 223.26, 225.86, 228.98, 230.59, 
    232.88, 232.64, 232.25, 241.4, 248.81, 257.52, 257.57, 255.79, 261.82, 
    267.65, 264.31, 254.1, 243.62, 232.08, 217.69, 205.14, 193.74,
  297.04, 296.74, 296.38, 295.92, 295.34, 294.69, 293.92, 293, 291.94, 
    290.74, 289.41, 287.98, 286.99, 285.1, 283.82, 291.75, 289.26, 287.34, 
    285.75, 283.69, 281.41, 279.28, 277.52, 276.21, 274.73, 272.94, 270.77, 
    269, 266.38, 263.31, 260.59, 257.3, 253.92, 250.1, 246.19, 242.71, 
    238.93, 235.01, 231.45, 228.44, 225.44, 222.29, 219.26, 216.09, 212.96, 
    209.59, 205.78, 202.2, 199.56, 197.58, 196.5, 196.76, 197.32, 197.74, 
    198.75, 199.73, 201.39, 204.27, 205.31, 208.75, 212.07, 211.66, 211.83, 
    212.58, 213.5, 216.18, 219.87, 222.58, 223.3, 222.46, 223.04, 226.2, 
    229.03, 230.06, 232.88, 232.93, 232.74, 241.22, 248.15, 257.72, 257.74, 
    255.95, 261.64, 267.77, 264.39, 254.07, 243.5, 232.06, 217.7, 205.25, 
    193.75,
  297.13, 296.83, 296.47, 296.01, 295.44, 294.79, 294.01, 293.1, 292.03, 
    290.83, 289.47, 288.01, 286.82, 285.15, 284.08, 291.59, 289.08, 287.35, 
    285.67, 283.61, 281.36, 279.28, 277.64, 276.32, 274.65, 272.85, 270.89, 
    269.13, 266.36, 263.27, 260.52, 257.26, 253.86, 250.09, 246.21, 242.72, 
    238.89, 235.01, 231.48, 228.36, 225.28, 222.2, 219.29, 216.11, 212.98, 
    209.68, 205.93, 202.34, 199.63, 197.55, 196.39, 196.54, 197.18, 198, 
    199.01, 199.8, 201.01, 204.02, 205.39, 208.81, 212.2, 211.81, 211.94, 
    212.66, 213.44, 215.99, 219.97, 222.63, 223.23, 222.38, 222.86, 226.47, 
    229.1, 229.63, 232.78, 233.11, 233.39, 241.06, 247.44, 257.81, 258.09, 
    256.03, 261.5, 267.75, 264.47, 254.09, 243.45, 232.04, 217.7, 205.28, 
    193.79,
  297.26, 296.96, 296.61, 296.15, 295.59, 294.93, 294.15, 293.24, 292.17, 
    290.96, 289.59, 288.09, 286.72, 285.18, 284.32, 291.41, 288.97, 287.37, 
    285.59, 283.51, 281.28, 279.29, 277.74, 276.33, 274.56, 272.83, 271.11, 
    269.26, 266.35, 263.26, 260.48, 257.24, 253.81, 250.08, 246.22, 242.7, 
    238.85, 235.01, 231.48, 228.27, 225.16, 222.14, 219.29, 216.1, 212.98, 
    209.75, 206.07, 202.48, 199.69, 197.54, 196.3, 196.29, 197, 198.26, 
    199.25, 199.92, 200.7, 203.71, 205.49, 208.85, 212.3, 211.97, 212.06, 
    212.74, 213.42, 215.79, 220.05, 222.64, 223.12, 222.34, 222.73, 226.62, 
    229.2, 229.36, 232.64, 233.18, 234.1, 240.89, 246.79, 257.79, 258.51, 
    256.09, 261.4, 267.71, 264.54, 254.13, 243.43, 232.01, 217.69, 205.28, 
    193.85,
  297.52, 297.24, 296.89, 296.44, 295.89, 295.25, 294.48, 293.6, 292.57, 
    291.36, 290, 288.37, 286.75, 285.26, 284.48, 290.55, 289.08, 287.42, 
    285.54, 283.42, 281.19, 279.29, 277.75, 276.19, 274.48, 272.86, 271.36, 
    269.38, 266.35, 263.27, 260.49, 257.26, 253.79, 250.07, 246.22, 242.63, 
    238.81, 235.01, 231.44, 228.18, 225.07, 222.14, 219.27, 216.07, 212.96, 
    209.8, 206.23, 202.63, 199.74, 197.51, 196.2, 196.03, 196.82, 198.54, 
    199.48, 200.01, 200.48, 203.41, 205.63, 208.84, 212.4, 212.13, 212.16, 
    212.75, 213.39, 215.69, 220.11, 222.63, 222.97, 222.32, 222.71, 226.72, 
    229.26, 229.17, 232.48, 233.17, 234.84, 240.8, 246.26, 257.59, 258.94, 
    256.15, 261.3, 267.61, 264.58, 254.23, 243.47, 231.98, 217.66, 205.23, 
    193.94,
  297.85, 297.58, 297.24, 296.8, 296.26, 295.62, 294.87, 294.01, 292.99, 
    291.78, 290.4, 288.65, 286.8, 285.25, 284.57, 289.84, 289.18, 287.42, 
    285.49, 283.35, 281.12, 279.32, 277.72, 276.03, 274.42, 272.9, 271.56, 
    269.46, 266.36, 263.29, 260.49, 257.28, 253.76, 250.07, 246.19, 242.53, 
    238.78, 235.02, 231.4, 228.09, 224.99, 222.16, 219.26, 216.04, 212.95, 
    209.85, 206.39, 202.77, 199.78, 197.49, 196.1, 195.76, 196.62, 198.81, 
    199.71, 200.11, 200.28, 203.13, 205.78, 208.83, 212.49, 212.3, 212.25, 
    212.75, 213.37, 215.6, 220.14, 222.64, 222.81, 222.31, 222.73, 226.77, 
    229.29, 229.04, 232.33, 233.12, 235.55, 240.72, 245.82, 257.35, 259.34, 
    256.21, 261.21, 267.51, 264.62, 254.33, 243.51, 231.94, 217.61, 205.16, 
    194.03,
  297.7, 297.44, 297.09, 296.63, 296.08, 295.44, 294.69, 293.81, 292.79, 
    291.63, 290.35, 288.93, 287.2, 285.71, 284.78, 288.34, 289.56, 287.39, 
    285.51, 283.37, 281.18, 279.36, 277.63, 275.94, 274.39, 272.96, 271.61, 
    269.44, 266.3, 263.25, 260.53, 257.31, 253.75, 250.06, 246.15, 242.47, 
    238.8, 235.05, 231.38, 228.02, 224.93, 222.16, 219.22, 216, 212.9, 
    209.87, 206.54, 202.94, 199.87, 197.51, 196.05, 195.46, 196.32, 198.94, 
    199.85, 200.13, 200.22, 203, 205.99, 208.87, 212.53, 212.47, 212.26, 
    212.64, 213.31, 215.66, 220.16, 222.62, 222.6, 222.27, 222.96, 226.74, 
    229.17, 229.03, 232.25, 233.03, 236.08, 240.66, 245.76, 256.91, 259.54, 
    256.34, 261.18, 267.36, 264.64, 254.48, 243.59, 231.89, 217.54, 205.05, 
    194.15,
  297.52, 297.26, 296.91, 296.45, 295.89, 295.24, 294.48, 293.59, 292.57, 
    291.44, 290.26, 289.16, 287.52, 286.26, 284.99, 286.82, 289.91, 287.37, 
    285.54, 283.41, 281.27, 279.39, 277.54, 275.92, 274.36, 273.02, 271.62, 
    269.39, 266.22, 263.18, 260.55, 257.34, 253.75, 250.05, 246.11, 242.43, 
    238.83, 235.09, 231.37, 227.95, 224.88, 222.15, 219.17, 215.94, 212.84, 
    209.88, 206.68, 203.12, 199.97, 197.58, 196.05, 195.17, 195.97, 198.98, 
    199.94, 200.12, 200.21, 202.96, 206.23, 208.99, 212.56, 212.61, 212.26, 
    212.49, 213.24, 215.72, 220.18, 222.62, 222.4, 222.22, 223.27, 226.66, 
    228.97, 229.05, 232.2, 233.01, 236.52, 240.54, 245.83, 256.46, 259.67, 
    256.48, 261.18, 267.21, 264.68, 254.61, 243.68, 231.82, 217.45, 204.94, 
    194.28,
  297.48, 297.2, 296.85, 296.39, 295.82, 295.16, 294.39, 293.49, 292.45, 
    291.31, 290.19, 289.25, 287.72, 286.86, 285.19, 285.87, 289.96, 287.33, 
    285.62, 283.49, 281.39, 279.41, 277.52, 275.97, 274.29, 273.12, 271.61, 
    269.28, 266.12, 263.14, 260.61, 257.37, 253.74, 250.03, 246.07, 242.43, 
    238.89, 235.12, 231.35, 227.88, 224.85, 222.14, 219.13, 215.88, 212.79, 
    209.87, 206.8, 203.28, 200.1, 197.75, 196.11, 194.91, 195.53, 198.85, 
    199.98, 200.11, 200.23, 203.02, 206.52, 209.18, 212.54, 212.75, 212.24, 
    212.28, 213.1, 215.81, 220.23, 222.62, 222.24, 222.17, 223.63, 226.57, 
    228.69, 229.09, 232.19, 233.02, 236.8, 240.4, 246.13, 256, 259.61, 
    256.71, 261.18, 267.06, 264.73, 254.77, 243.77, 231.74, 217.33, 204.84, 
    194.41,
  297.52, 297.22, 296.85, 296.4, 295.83, 295.17, 294.4, 293.48, 292.43, 
    291.27, 290.21, 289.32, 287.83, 287.35, 285.35, 285.09, 289.94, 287.32, 
    285.72, 283.57, 281.49, 279.4, 277.53, 276.04, 274.21, 273.21, 271.58, 
    269.14, 266.01, 263.12, 260.67, 257.39, 253.73, 250, 246.04, 242.45, 
    238.95, 235.16, 231.32, 227.81, 224.82, 222.14, 219.1, 215.83, 212.74, 
    209.86, 206.9, 203.42, 200.23, 197.95, 196.21, 194.68, 195.04, 198.64, 
    200, 200.11, 200.27, 203.1, 206.83, 209.41, 212.52, 212.87, 212.24, 
    212.03, 212.93, 215.9, 220.29, 222.64, 222.1, 222.11, 224, 226.48, 
    228.37, 229.14, 232.17, 233.09, 237.02, 240.2, 246.48, 255.55, 259.51, 
    256.97, 261.17, 266.92, 264.79, 254.92, 243.86, 231.66, 217.2, 204.75, 
    194.53,
  297.58, 297.3, 296.95, 296.5, 295.94, 295.28, 294.51, 293.6, 292.56, 
    291.43, 290.38, 289.35, 287.91, 287.37, 285.43, 284.66, 289.55, 287.36, 
    285.85, 283.62, 281.43, 279.32, 277.51, 276.05, 274.18, 273.2, 271.54, 
    268.96, 265.87, 263.17, 260.74, 257.39, 253.69, 249.93, 246.03, 242.5, 
    238.99, 235.15, 231.27, 227.74, 224.78, 222.13, 219.1, 215.76, 212.66, 
    209.86, 206.99, 203.56, 200.4, 198.18, 196.29, 194.53, 194.51, 198.29, 
    199.95, 200.07, 200.34, 203.35, 207.22, 209.72, 212.41, 212.89, 212.19, 
    211.77, 212.72, 216.08, 220.43, 222.59, 221.95, 222.07, 224.37, 226.43, 
    228, 229.11, 232.15, 233.35, 237.19, 239.94, 246.72, 255.25, 259.26, 
    257.33, 261.11, 266.87, 264.86, 255.07, 243.9, 231.57, 217.03, 204.71, 
    194.62,
  297.64, 297.38, 297.05, 296.6, 296.04, 295.38, 294.62, 293.71, 292.67, 
    291.55, 290.49, 289.4, 287.96, 287.28, 285.57, 284.49, 289.14, 287.39, 
    285.97, 283.67, 281.34, 279.23, 277.47, 276.05, 274.18, 273.12, 271.49, 
    268.78, 265.72, 263.27, 260.82, 257.38, 253.64, 249.84, 246.02, 242.56, 
    239.03, 235.13, 231.23, 227.68, 224.76, 222.12, 219.08, 215.67, 212.57, 
    209.86, 207.09, 203.71, 200.58, 198.42, 196.36, 194.4, 193.95, 197.91, 
    199.89, 200.04, 200.38, 203.6, 207.62, 210.04, 212.3, 212.87, 212.14, 
    211.53, 212.52, 216.27, 220.57, 222.55, 221.83, 222.03, 224.69, 226.43, 
    227.67, 229.02, 232.09, 233.65, 237.36, 239.67, 246.89, 255, 258.97, 
    257.74, 261.01, 266.86, 264.92, 255.23, 243.91, 231.49, 216.85, 204.71, 
    194.69,
  297.62, 297.36, 297.03, 296.58, 296.02, 295.36, 294.59, 293.69, 292.66, 
    291.53, 290.53, 289.39, 288.05, 287.27, 285.73, 284.6, 288.95, 287.38, 
    286.03, 283.72, 281.32, 279.16, 277.39, 276.04, 274.21, 272.97, 271.42, 
    268.64, 265.62, 263.41, 260.9, 257.37, 253.58, 249.76, 246.04, 242.62, 
    239.04, 235.11, 231.19, 227.64, 224.75, 222.12, 219.06, 215.58, 212.5, 
    209.87, 207.18, 203.87, 200.75, 198.61, 196.44, 194.3, 193.42, 197.56, 
    199.84, 200.01, 200.4, 203.83, 208.02, 210.36, 212.17, 212.8, 212.1, 
    211.33, 212.36, 216.44, 220.68, 222.5, 221.73, 221.98, 224.94, 226.5, 
    227.42, 228.85, 231.96, 233.98, 237.55, 239.44, 246.98, 254.81, 258.62, 
    258.18, 260.89, 266.9, 265, 255.37, 243.89, 231.41, 216.67, 204.75, 194.75,
  297.51, 297.26, 296.91, 296.45, 295.9, 295.24, 294.47, 293.56, 292.55, 
    291.41, 290.54, 289.32, 288.13, 287.34, 285.9, 284.85, 288.85, 287.33, 
    286.03, 283.79, 281.34, 279.1, 277.29, 276.03, 274.27, 272.79, 271.3, 
    268.51, 265.56, 263.58, 260.95, 257.34, 253.52, 249.68, 246.06, 242.68, 
    239.04, 235.09, 231.15, 227.61, 224.76, 222.13, 219.03, 215.51, 212.46, 
    209.88, 207.25, 204.04, 200.92, 198.77, 196.51, 194.21, 192.91, 197.24, 
    199.8, 199.98, 200.4, 204.04, 208.39, 210.66, 212.04, 212.67, 212.07, 
    211.2, 212.25, 216.61, 220.74, 222.43, 221.66, 221.95, 225.1, 226.65, 
    227.26, 228.61, 231.8, 234.32, 237.74, 239.28, 246.99, 254.65, 258.24, 
    258.63, 260.75, 266.98, 265.07, 255.5, 243.83, 231.32, 216.49, 204.82, 
    194.78,
  297.4, 297.13, 296.78, 296.33, 295.77, 295.11, 294.35, 293.44, 292.41, 
    291.39, 290.54, 289.31, 288.28, 287.55, 286.01, 284.96, 288.8, 287.26, 
    286, 283.84, 281.36, 279.02, 277.22, 276.09, 274.36, 272.64, 271.06, 
    268.34, 265.6, 263.76, 260.98, 257.29, 253.45, 249.65, 246.11, 242.75, 
    239.03, 235.05, 231.11, 227.62, 224.78, 222.15, 219, 215.48, 212.47, 
    209.91, 207.3, 204.19, 201.1, 198.87, 196.55, 194.11, 192.47, 196.96, 
    199.8, 199.96, 200.37, 204.16, 208.65, 210.89, 211.89, 212.5, 212.08, 
    211.2, 212.26, 216.74, 220.71, 222.27, 221.62, 222, 225.17, 226.87, 
    227.21, 228.27, 231.65, 234.62, 237.81, 239.28, 246.95, 254.54, 257.86, 
    259.01, 260.6, 267.2, 265.12, 255.6, 243.7, 231.26, 216.33, 204.94, 194.78,
  297.3, 297.04, 296.7, 296.25, 295.7, 295.04, 294.27, 293.37, 292.3, 291.48, 
    290.55, 289.41, 288.45, 287.8, 286.08, 285, 288.73, 287.21, 286.02, 
    283.88, 281.38, 278.96, 277.22, 276.19, 274.46, 272.5, 270.76, 268.15, 
    265.69, 263.92, 261, 257.23, 253.38, 249.64, 246.18, 242.82, 239, 235.01, 
    231.09, 227.66, 224.83, 222.18, 218.97, 215.45, 212.5, 209.95, 207.33, 
    204.32, 201.29, 198.95, 196.59, 194.01, 192.09, 196.68, 199.82, 199.95, 
    200.35, 204.18, 208.83, 211.11, 211.76, 212.31, 212.1, 211.26, 212.35, 
    216.83, 220.62, 222.1, 221.61, 222.07, 225.24, 227.12, 227.2, 227.91, 
    231.46, 234.92, 237.81, 239.33, 246.95, 254.47, 257.46, 259.29, 260.48, 
    267.48, 265.17, 255.67, 243.53, 231.2, 216.19, 205.07, 194.77,
  297.16, 296.89, 296.56, 296.12, 295.57, 294.92, 294.15, 293.26, 292.2, 
    291.51, 290.54, 289.58, 288.61, 287.98, 286.2, 285.02, 288.47, 287.19, 
    286.08, 283.94, 281.43, 278.97, 277.29, 276.32, 274.55, 272.35, 270.44, 
    267.98, 265.8, 264.07, 261.01, 257.17, 253.31, 249.66, 246.24, 242.86, 
    238.96, 234.96, 231.08, 227.71, 224.89, 222.21, 218.93, 215.41, 212.53, 
    210, 207.37, 204.42, 201.46, 199.03, 196.62, 193.9, 191.79, 196.38, 
    199.88, 199.97, 200.35, 204.13, 208.96, 211.33, 211.66, 212.11, 212.11, 
    211.35, 212.51, 216.88, 220.48, 221.91, 221.6, 222.15, 225.32, 227.36, 
    227.2, 227.57, 231.26, 235.2, 237.75, 239.41, 246.99, 254.43, 257.05, 
    259.47, 260.44, 267.8, 265.19, 255.69, 243.34, 231.16, 216.09, 205.21, 
    194.76,
  296.89, 296.62, 296.28, 295.83, 295.27, 294.63, 293.88, 293.01, 292.14, 
    291.4, 290.5, 289.75, 288.72, 288.03, 286.36, 284.98, 287.81, 287.11, 
    286.11, 284, 281.52, 279.05, 277.42, 276.39, 274.56, 272.17, 270.11, 
    267.83, 265.92, 264.17, 261, 257.09, 253.26, 249.73, 246.32, 242.84, 
    238.9, 234.92, 231.11, 227.75, 224.93, 222.22, 218.86, 215.36, 212.56, 
    210.08, 207.42, 204.49, 201.59, 199.11, 196.62, 193.8, 191.6, 196.03, 
    199.98, 200.02, 200.44, 204.04, 208.97, 211.49, 211.62, 211.9, 212.12, 
    211.47, 212.69, 216.9, 220.3, 221.71, 221.64, 222.27, 225.41, 227.55, 
    227.22, 227.28, 231.07, 235.39, 237.62, 239.52, 247.17, 254.38, 256.68, 
    259.41, 260.59, 268.15, 265.17, 255.61, 243.15, 231.12, 216.05, 205.31, 
    194.78,
  296.64, 296.36, 296, 295.55, 294.98, 294.36, 293.62, 292.77, 292.11, 
    291.32, 290.52, 289.89, 288.83, 288.05, 286.49, 285.02, 287.16, 286.91, 
    286.05, 284.06, 281.63, 279.17, 277.54, 276.43, 274.54, 272.01, 269.84, 
    267.73, 266.04, 264.23, 260.97, 257.02, 253.22, 249.81, 246.4, 242.81, 
    238.85, 234.9, 231.16, 227.8, 224.96, 222.21, 218.78, 215.29, 212.57, 
    210.17, 207.5, 204.55, 201.67, 199.15, 196.6, 193.68, 191.45, 195.67, 
    200.09, 200.11, 200.6, 203.97, 208.93, 211.6, 211.63, 211.7, 212.09, 
    211.58, 212.88, 216.9, 220.13, 221.53, 221.73, 222.4, 225.48, 227.67, 
    227.26, 227.06, 230.91, 235.49, 237.46, 239.66, 247.45, 254.27, 256.37, 
    259.21, 260.93, 268.44, 265.15, 255.46, 242.99, 231.08, 216.07, 205.37, 
    194.82,
  296.41, 296.12, 295.77, 295.33, 294.78, 294.15, 293.44, 292.61, 292.16, 
    291.31, 290.65, 290, 288.99, 288.1, 286.67, 285.23, 286.38, 286.68, 
    285.98, 284.14, 281.76, 279.31, 277.63, 276.47, 274.57, 271.94, 269.69, 
    267.7, 266.16, 264.26, 260.93, 256.97, 253.24, 249.91, 246.48, 242.76, 
    238.83, 234.92, 231.23, 227.87, 225, 222.2, 218.69, 215.19, 212.53, 
    210.25, 207.61, 204.63, 201.72, 199.13, 196.55, 193.55, 191.36, 195.38, 
    200.14, 200.23, 200.78, 203.93, 208.88, 211.69, 211.68, 211.52, 212.02, 
    211.65, 213.09, 216.9, 219.97, 221.38, 221.8, 222.54, 225.53, 227.69, 
    227.3, 226.95, 230.78, 235.51, 237.25, 239.79, 247.79, 254.15, 256.11, 
    258.92, 261.46, 268.63, 265.07, 255.22, 242.86, 231.06, 216.15, 205.38, 
    194.88,
  296.18, 295.9, 295.56, 295.11, 294.58, 293.96, 293.25, 292.49, 292.2, 
    291.31, 290.79, 290.13, 289.16, 288.21, 286.9, 285.5, 285.51, 286.4, 
    285.91, 284.24, 281.91, 279.46, 277.7, 276.52, 274.6, 271.9, 269.58, 
    267.71, 266.28, 264.28, 260.89, 256.92, 253.25, 250, 246.56, 242.73, 
    238.82, 234.96, 231.31, 227.95, 225.05, 222.18, 218.61, 215.08, 212.46, 
    210.32, 207.74, 204.72, 201.76, 199.11, 196.49, 193.41, 191.24, 195.11, 
    200.17, 200.38, 200.99, 203.88, 208.84, 211.77, 211.75, 211.34, 211.91, 
    211.72, 213.32, 216.92, 219.82, 221.26, 221.87, 222.67, 225.54, 227.68, 
    227.33, 226.92, 230.66, 235.49, 237.03, 239.93, 248.14, 254, 255.88, 
    258.61, 262.08, 268.73, 265, 254.96, 242.77, 231.04, 216.26, 205.37, 
    194.95,
  296.25, 295.97, 295.62, 295.19, 294.67, 294.05, 293.33, 292.64, 292.21, 
    291.38, 290.77, 290.1, 289.18, 288.21, 287, 285.58, 285, 286.03, 285.81, 
    284.24, 281.96, 279.53, 277.71, 276.55, 274.59, 271.86, 269.56, 267.8, 
    266.39, 264.25, 260.81, 256.87, 253.26, 250.03, 246.57, 242.7, 238.82, 
    235.02, 231.38, 228.02, 225.1, 222.14, 218.51, 214.95, 212.33, 210.3, 
    207.86, 204.85, 201.81, 199.05, 196.39, 193.22, 191.14, 194.94, 200.09, 
    200.55, 201.14, 203.96, 208.84, 211.82, 211.87, 211.29, 211.83, 211.69, 
    213.47, 216.93, 219.7, 221.2, 221.91, 222.85, 225.5, 227.5, 227.31, 
    227.15, 230.6, 235.34, 236.79, 240.09, 248.54, 253.81, 255.69, 258.39, 
    262.89, 268.53, 264.91, 254.63, 242.8, 231.01, 216.41, 205.3, 195.06,
  296.2, 295.92, 295.57, 295.15, 294.63, 294, 293.29, 292.7, 292.17, 291.42, 
    290.77, 290.08, 289.22, 288.25, 287.19, 285.72, 284.46, 285.48, 285.63, 
    284.18, 281.98, 279.58, 277.75, 276.61, 274.58, 271.83, 269.57, 267.92, 
    266.5, 264.2, 260.71, 256.8, 253.25, 250.05, 246.56, 242.67, 238.83, 
    235.07, 231.45, 228.08, 225.15, 222.1, 218.41, 214.83, 212.21, 210.27, 
    207.96, 204.97, 201.87, 199, 196.28, 193.06, 191.02, 194.76, 200, 200.72, 
    201.28, 204.03, 208.86, 211.87, 211.99, 211.3, 211.76, 211.64, 213.57, 
    216.91, 219.61, 221.18, 221.95, 223.01, 225.44, 227.33, 227.26, 227.43, 
    230.55, 235.19, 236.53, 240.25, 248.92, 253.63, 255.5, 258.22, 263.7, 
    268.23, 264.82, 254.31, 242.86, 230.98, 216.57, 205.21, 195.17,
  296.11, 295.83, 295.49, 295.06, 294.53, 293.91, 293.18, 292.61, 292, 
    291.32, 290.75, 290.05, 289.27, 288.33, 287.32, 285.82, 284.49, 284.83, 
    285.42, 284.1, 281.99, 279.65, 277.84, 276.65, 274.55, 271.84, 269.63, 
    268.07, 266.61, 264.18, 260.64, 256.76, 253.26, 250.06, 246.54, 242.68, 
    238.86, 235.14, 231.52, 228.16, 225.22, 222.08, 218.33, 214.73, 212.1, 
    210.18, 207.98, 205.1, 201.96, 198.97, 196.18, 192.93, 190.83, 194.55, 
    199.95, 200.89, 201.36, 204.15, 208.86, 211.97, 212.16, 211.35, 211.7, 
    211.55, 213.62, 216.86, 219.55, 221.2, 221.99, 223.15, 225.38, 227.13, 
    227.17, 227.72, 230.57, 235.07, 236.3, 240.38, 249.16, 253.48, 255.46, 
    258.18, 264.4, 267.78, 264.72, 254.04, 242.97, 230.97, 216.71, 205.11, 
    195.27,
  296.03, 295.74, 295.4, 294.98, 294.44, 293.81, 293.05, 292.48, 291.77, 
    291.23, 290.73, 290.02, 289.31, 288.41, 287.44, 286.03, 284.57, 284.14, 
    285.21, 284.03, 282, 279.72, 277.95, 276.69, 274.54, 271.87, 269.69, 
    268.23, 266.73, 264.17, 260.57, 256.71, 253.27, 250.07, 246.54, 242.68, 
    238.89, 235.21, 231.6, 228.25, 225.28, 222.07, 218.25, 214.64, 212.01, 
    210.09, 207.99, 205.21, 202.07, 198.96, 196.09, 192.82, 190.64, 194.34, 
    199.92, 201.04, 201.44, 204.23, 208.83, 212.09, 212.36, 211.44, 211.65, 
    211.45, 213.63, 216.78, 219.5, 221.26, 222.01, 223.26, 225.34, 226.97, 
    227.03, 228, 230.61, 234.96, 236.09, 240.5, 249.34, 253.35, 255.47, 
    258.18, 265.03, 267.29, 264.62, 253.8, 243.1, 230.96, 216.84, 205.02, 
    195.36,
  296.06, 295.78, 295.45, 295.02, 294.48, 293.84, 293.11, 292.54, 291.74, 
    291.26, 290.71, 290.04, 289.35, 288.45, 287.39, 286.01, 284.69, 284.13, 
    284.94, 283.85, 281.94, 279.73, 277.96, 276.64, 274.49, 271.9, 269.77, 
    268.36, 266.83, 264.17, 260.52, 256.69, 253.28, 250.05, 246.52, 242.66, 
    238.91, 235.26, 231.66, 228.32, 225.32, 222.05, 218.19, 214.55, 211.92, 
    209.98, 207.95, 205.33, 202.21, 199, 196.02, 192.73, 190.46, 194.1, 
    199.96, 201.17, 201.61, 204.27, 208.62, 212.21, 212.6, 211.62, 211.67, 
    211.34, 213.52, 216.59, 219.54, 221.39, 222, 223.35, 225.4, 226.82, 
    226.76, 228.24, 230.74, 234.9, 235.96, 240.57, 249.3, 253.32, 255.67, 
    258.24, 265.33, 266.81, 264.55, 253.68, 243.24, 230.96, 216.92, 204.96, 
    195.43,
  296.1, 295.83, 295.5, 295.07, 294.54, 293.89, 293.19, 292.63, 291.73, 
    291.29, 290.68, 290.04, 289.37, 288.47, 287.33, 285.94, 284.74, 284.24, 
    284.69, 283.67, 281.87, 279.73, 277.99, 276.6, 274.44, 271.92, 269.82, 
    268.44, 266.91, 264.17, 260.48, 256.67, 253.29, 250.03, 246.5, 242.65, 
    238.91, 235.31, 231.72, 228.39, 225.34, 222.02, 218.14, 214.45, 211.82, 
    209.87, 207.91, 205.44, 202.36, 199.07, 195.96, 192.65, 190.29, 193.87, 
    200.01, 201.3, 201.79, 204.28, 208.39, 212.31, 212.84, 211.8, 211.68, 
    211.23, 213.4, 216.38, 219.59, 221.55, 222, 223.41, 225.5, 226.67, 
    226.45, 228.47, 230.87, 234.87, 235.85, 240.65, 249.14, 253.32, 255.94, 
    258.33, 265.49, 266.38, 264.49, 253.6, 243.36, 230.97, 216.98, 204.91, 
    195.48,
  296.12, 295.85, 295.53, 295.1, 294.57, 293.93, 293.25, 292.81, 291.89, 
    291.32, 290.71, 290.03, 289.38, 288.47, 287.31, 285.89, 284.71, 284.46, 
    284.56, 283.54, 281.84, 279.74, 278.01, 276.56, 274.39, 271.93, 269.84, 
    268.48, 266.93, 264.14, 260.43, 256.66, 253.33, 250.03, 246.49, 242.65, 
    238.93, 235.34, 231.78, 228.47, 225.38, 222, 218.09, 214.36, 211.69, 
    209.75, 207.85, 205.53, 202.51, 199.15, 195.92, 192.59, 190.14, 193.69, 
    200.08, 201.45, 202.01, 204.22, 208.18, 212.33, 213.07, 212.01, 211.68, 
    211.11, 213.23, 216.16, 219.69, 221.77, 222.03, 223.46, 225.6, 226.46, 
    226.15, 228.69, 231.02, 234.86, 235.76, 240.77, 248.81, 253.38, 256.33, 
    258.44, 265.37, 266.08, 264.45, 253.59, 243.46, 231.01, 216.98, 204.9, 
    195.5,
  296.15, 295.88, 295.56, 295.13, 294.6, 293.97, 293.31, 292.98, 292.15, 
    291.38, 290.79, 290.07, 289.38, 288.47, 287.34, 285.93, 284.64, 284.69, 
    284.57, 283.49, 281.84, 279.78, 278.06, 276.55, 274.37, 271.94, 269.82, 
    268.46, 266.9, 264.1, 260.38, 256.66, 253.39, 250.05, 246.48, 242.66, 
    238.96, 235.39, 231.87, 228.56, 225.43, 221.97, 218.05, 214.29, 211.53, 
    209.57, 207.79, 205.61, 202.66, 199.26, 195.91, 192.56, 190.06, 193.57, 
    200.12, 201.6, 202.22, 204.14, 207.97, 212.31, 213.27, 212.19, 211.67, 
    211.01, 213.05, 215.95, 219.82, 221.98, 222.1, 223.54, 225.69, 226.17, 
    225.92, 228.89, 231.13, 234.85, 235.74, 240.98, 248.28, 253.49, 256.78, 
    258.56, 265.02, 265.96, 264.39, 253.66, 243.51, 231.06, 216.94, 204.92, 
    195.5,
  296.25, 295.99, 295.65, 295.22, 294.69, 294.07, 293.42, 293.02, 292.3, 
    291.45, 290.81, 290.08, 289.34, 288.43, 287.38, 286.05, 284.62, 284.91, 
    284.59, 283.47, 281.88, 279.86, 278.11, 276.54, 274.35, 271.94, 269.8, 
    268.38, 266.82, 264.01, 260.32, 256.66, 253.45, 250.09, 246.48, 242.66, 
    238.99, 235.44, 231.96, 228.66, 225.46, 221.94, 218.01, 214.25, 211.34, 
    209.31, 207.73, 205.69, 202.79, 199.36, 195.93, 192.54, 190.09, 193.54, 
    200.08, 201.77, 202.38, 204.08, 207.8, 212.25, 213.43, 212.33, 211.64, 
    210.91, 212.86, 215.79, 220, 222.17, 222.19, 223.62, 225.7, 225.82, 
    225.85, 229.04, 231.18, 234.76, 235.83, 241.29, 247.58, 253.65, 257.25, 
    258.69, 264.45, 266.07, 264.3, 253.81, 243.51, 231.14, 216.85, 204.99, 
    195.47,
  296.34, 296.07, 295.72, 295.28, 294.76, 294.16, 293.51, 292.98, 292.35, 
    291.49, 290.77, 290.05, 289.26, 288.37, 287.43, 286.16, 284.61, 285.08, 
    284.57, 283.45, 281.93, 279.93, 278.15, 276.52, 274.31, 271.93, 269.77, 
    268.29, 266.73, 263.89, 260.23, 256.66, 253.51, 250.11, 246.46, 242.65, 
    239, 235.5, 232.07, 228.76, 225.47, 221.9, 217.98, 214.21, 211.15, 
    209.01, 207.68, 205.78, 202.89, 199.43, 195.96, 192.53, 190.19, 193.54, 
    199.99, 201.97, 202.5, 204.05, 207.71, 212.17, 213.56, 212.44, 211.56, 
    210.78, 212.69, 215.7, 220.21, 222.34, 222.29, 223.69, 225.66, 225.45, 
    225.85, 229.16, 231.26, 234.62, 235.99, 241.64, 246.81, 253.83, 257.69, 
    258.8, 263.8, 266.31, 264.2, 253.99, 243.48, 231.22, 216.73, 205.07, 
    195.43 ;

 temp_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 shum =
  0.011025, 0.010689, 0.01055, 0.010469, 0.010416, 0.010376, 0.010344, 
    0.010319, 0.010301, 0.01028, 0.010242, 0.010062, 0.0091736, 0.0090951, 
    0.0088283, 0.0012647, 0.0012706, 0.001471, 0.0012792, 0.0012191, 
    0.001081, 0.00077981, 0.00047109, 0.00025036, 0.00016494, 0.000141, 
    0.00014109, 0.0001252, 9.4174e-05, 0.00013455, 0.00055901, 0.0005074, 
    0.00027088, 0.00025257, 0.00024511, 0.00016537, 0.00012688, 0.00011139, 
    8.5684e-05, 5.2974e-05, 3.0922e-05, 2.0495e-05, 1.795e-05, 1.5492e-05, 
    1.1227e-05, 1.2245e-05, 1.5283e-05, 9.7364e-06, 6.35e-06, 4.7917e-06, 
    4.4182e-06, 3.9087e-06, 3.6979e-06, 3.5102e-06, 3.1083e-06, 2.8547e-06, 
    2.6855e-06, 2.5881e-06, 2.5498e-06, 2.4835e-06, 2.4448e-06, 2.4449e-06, 
    2.4651e-06, 2.4966e-06, 2.5491e-06, 2.6167e-06, 2.6957e-06, 2.7599e-06, 
    2.7972e-06, 2.8235e-06, 2.8408e-06, 2.847e-06, 2.8484e-06, 2.8621e-06, 
    2.9096e-06, 2.9778e-06, 3.0633e-06, 3.2255e-06, 3.397e-06, 3.587e-06, 
    3.6608e-06, 3.6367e-06, 3.6985e-06, 3.9468e-06, 3.9485e-06, 3.8956e-06, 
    3.9625e-06, 4.0027e-06, 3.9995e-06, 3.8839e-06, 2.6092e-06,
  0.011086, 0.010755, 0.010618, 0.010538, 0.010486, 0.010446, 0.010414, 
    0.01039, 0.010372, 0.010352, 0.010314, 0.010117, 0.0091823, 0.0090461, 
    0.0085294, 0.0011735, 0.0011907, 0.0014253, 0.0012745, 0.0011734, 
    0.0010458, 0.00078516, 0.00046486, 0.00024143, 0.00020532, 0.00015646, 
    0.000149, 0.00012279, 8.7212e-05, 0.00013971, 0.0006278, 0.00055679, 
    0.00028794, 0.00024431, 0.00024014, 0.00015665, 0.00012712, 0.00011314, 
    8.3374e-05, 5.117e-05, 3.1091e-05, 2.1999e-05, 1.9361e-05, 1.6919e-05, 
    1.2052e-05, 1.1425e-05, 1.5449e-05, 9.8346e-06, 6.3206e-06, 4.8451e-06, 
    4.4651e-06, 3.8939e-06, 3.6132e-06, 3.4732e-06, 3.1056e-06, 2.8464e-06, 
    2.6886e-06, 2.5858e-06, 2.5451e-06, 2.4818e-06, 2.4449e-06, 2.4451e-06, 
    2.4649e-06, 2.4971e-06, 2.5487e-06, 2.6146e-06, 2.6947e-06, 2.7602e-06, 
    2.7968e-06, 2.8233e-06, 2.8406e-06, 2.8465e-06, 2.8477e-06, 2.8607e-06, 
    2.9087e-06, 2.9794e-06, 3.0654e-06, 3.2235e-06, 3.3934e-06, 3.5854e-06, 
    3.6573e-06, 3.6344e-06, 3.6907e-06, 3.9443e-06, 3.9468e-06, 3.8947e-06, 
    3.9633e-06, 4.0032e-06, 3.9999e-06, 3.8782e-06, 2.6136e-06,
  0.011141, 0.010812, 0.010676, 0.010596, 0.010543, 0.010503, 0.010472, 
    0.010448, 0.010432, 0.010416, 0.010383, 0.010185, 0.0093977, 0.009234, 
    0.0082472, 0.0010907, 0.0011556, 0.0013756, 0.0012962, 0.0011678, 
    0.001025, 0.00076992, 0.00044523, 0.0002741, 0.0002739, 0.00017311, 
    0.00015258, 0.00011233, 8.0453e-05, 0.00016152, 0.00065549, 0.00059149, 
    0.00031455, 0.0002385, 0.00023497, 0.00015401, 0.00013233, 0.00011126, 
    7.869e-05, 4.9492e-05, 3.1329e-05, 2.3279e-05, 2.0284e-05, 1.7931e-05, 
    1.2914e-05, 1.0766e-05, 1.5038e-05, 9.7986e-06, 6.3828e-06, 4.8808e-06, 
    4.4655e-06, 3.8978e-06, 3.5174e-06, 3.4259e-06, 3.1038e-06, 2.8371e-06, 
    2.6905e-06, 2.5852e-06, 2.539e-06, 2.4802e-06, 2.4447e-06, 2.4454e-06, 
    2.465e-06, 2.4973e-06, 2.5483e-06, 2.6119e-06, 2.694e-06, 2.7593e-06, 
    2.7966e-06, 2.8234e-06, 2.8404e-06, 2.846e-06, 2.8472e-06, 2.8591e-06, 
    2.9074e-06, 2.9797e-06, 3.0695e-06, 3.2221e-06, 3.3902e-06, 3.5819e-06, 
    3.6481e-06, 3.6287e-06, 3.6877e-06, 3.9412e-06, 3.9458e-06, 3.8937e-06, 
    3.9643e-06, 4.0034e-06, 4.0001e-06, 3.8747e-06, 2.6162e-06,
  0.011131, 0.010803, 0.010666, 0.010585, 0.01053, 0.010489, 0.010454, 
    0.010423, 0.010403, 0.010389, 0.010342, 0.010149, 0.0095515, 0.0094059, 
    0.0083193, 0.0010615, 0.0011268, 0.0013334, 0.0013179, 0.0011851, 
    0.0010216, 0.00075285, 0.00043931, 0.00034469, 0.00036142, 0.00018826, 
    0.00015038, 9.8835e-05, 7.6226e-05, 0.00018839, 0.00068154, 0.00062385, 
    0.00034496, 0.00023649, 0.00023076, 0.00015599, 0.00013588, 0.00010744, 
    7.4326e-05, 4.8267e-05, 3.1553e-05, 2.4152e-05, 2.0817e-05, 1.8384e-05, 
    1.3445e-05, 1.0317e-05, 1.4152e-05, 9.9588e-06, 6.5024e-06, 4.9298e-06, 
    4.4815e-06, 3.9208e-06, 3.4346e-06, 3.3786e-06, 3.1032e-06, 2.8248e-06, 
    2.6909e-06, 2.5852e-06, 2.5329e-06, 2.4789e-06, 2.4441e-06, 2.4457e-06, 
    2.4652e-06, 2.4975e-06, 2.5481e-06, 2.6093e-06, 2.6936e-06, 2.7579e-06, 
    2.796e-06, 2.8235e-06, 2.8403e-06, 2.8455e-06, 2.8467e-06, 2.858e-06, 
    2.9061e-06, 2.979e-06, 3.0746e-06, 3.2205e-06, 3.3872e-06, 3.5771e-06, 
    3.6353e-06, 3.6207e-06, 3.6862e-06, 3.9381e-06, 3.945e-06, 3.8925e-06, 
    3.9657e-06, 4.0034e-06, 4.0002e-06, 3.8701e-06, 2.616e-06,
  0.011075, 0.010728, 0.01058, 0.01049, 0.010425, 0.010374, 0.010317, 
    0.010246, 0.0102, 0.010191, 0.010141, 0.010057, 0.0097793, 0.0096411, 
    0.0087785, 0.0013293, 0.0011155, 0.001291, 0.0013248, 0.001224, 
    0.0010421, 0.00075226, 0.00047637, 0.00046927, 0.00047312, 0.00021363, 
    0.00014109, 8.4649e-05, 7.3012e-05, 0.0002235, 0.00071805, 0.00064524, 
    0.00036791, 0.0002386, 0.00022993, 0.00016506, 0.00013485, 0.00010132, 
    7.1942e-05, 4.7181e-05, 3.171e-05, 2.4339e-05, 2.0861e-05, 1.8241e-05, 
    1.3621e-05, 1.033e-05, 1.2624e-05, 1.0386e-05, 6.7126e-06, 5.0134e-06, 
    4.5387e-06, 3.9647e-06, 3.3803e-06, 3.3424e-06, 3.0973e-06, 2.8218e-06, 
    2.6908e-06, 2.5858e-06, 2.5266e-06, 2.4776e-06, 2.4434e-06, 2.4459e-06, 
    2.4654e-06, 2.4975e-06, 2.5474e-06, 2.6068e-06, 2.6932e-06, 2.7566e-06, 
    2.7956e-06, 2.8237e-06, 2.8402e-06, 2.845e-06, 2.8462e-06, 2.8574e-06, 
    2.905e-06, 2.9783e-06, 3.08e-06, 3.2201e-06, 3.3845e-06, 3.5714e-06, 
    3.6172e-06, 3.6065e-06, 3.6825e-06, 3.9359e-06, 3.9448e-06, 3.8911e-06, 
    3.9672e-06, 4.0035e-06, 4.0003e-06, 3.8631e-06, 2.6136e-06,
  0.01091, 0.010542, 0.010383, 0.010286, 0.010216, 0.01016, 0.010107, 
    0.010051, 0.010014, 0.0099891, 0.0099198, 0.0098762, 0.0099197, 
    0.0098195, 0.008861, 0.0014808, 0.0010831, 0.0012403, 0.0013274, 
    0.0012609, 0.0010601, 0.00074806, 0.00053222, 0.00061528, 0.00058993, 
    0.00024242, 0.00013097, 7.1791e-05, 6.995e-05, 0.0002626, 0.00075886, 
    0.00066817, 0.0003923, 0.00024156, 0.0002318, 0.0001754, 0.00013279, 
    9.4483e-05, 6.9687e-05, 4.5779e-05, 3.1768e-05, 2.4292e-05, 2.0706e-05, 
    1.7845e-05, 1.3579e-05, 1.0469e-05, 1.0967e-05, 1.0764e-05, 6.9408e-06, 
    5.1048e-06, 4.6127e-06, 4.0286e-06, 3.339e-06, 3.3078e-06, 3.0917e-06, 
    2.8194e-06, 2.6904e-06, 2.5869e-06, 2.5216e-06, 2.4769e-06, 2.4428e-06, 
    2.4462e-06, 2.4656e-06, 2.4974e-06, 2.5469e-06, 2.6044e-06, 2.6926e-06, 
    2.7552e-06, 2.795e-06, 2.824e-06, 2.8403e-06, 2.8446e-06, 2.8457e-06, 
    2.8572e-06, 2.904e-06, 2.978e-06, 3.0853e-06, 3.2197e-06, 3.3819e-06, 
    3.5656e-06, 3.5978e-06, 3.59e-06, 3.6779e-06, 3.9343e-06, 3.9446e-06, 
    3.8896e-06, 3.9689e-06, 4.0035e-06, 4.0004e-06, 3.8546e-06, 2.6101e-06,
  0.011287, 0.010943, 0.010796, 0.010707, 0.010642, 0.010587, 0.01053, 
    0.010434, 0.01033, 0.010208, 0.010034, 0.0099479, 0.0099216, 0.0098003, 
    0.0088584, 0.0026757, 0.0010383, 0.0011423, 0.001329, 0.0013017, 
    0.0010775, 0.00077795, 0.00066542, 0.00083789, 0.00088118, 0.00026364, 
    0.00011784, 6.1784e-05, 9.6857e-05, 0.00037592, 0.00079783, 0.0006776, 
    0.00040637, 0.00025051, 0.00024119, 0.00017998, 0.00012561, 8.9313e-05, 
    6.7916e-05, 4.4978e-05, 3.1846e-05, 2.3975e-05, 1.9812e-05, 1.6785e-05, 
    1.3223e-05, 1.0662e-05, 9.9202e-06, 1.0608e-05, 7.1413e-06, 5.2383e-06, 
    4.7605e-06, 4.1083e-06, 3.3075e-06, 3.2771e-06, 3.0863e-06, 2.8196e-06, 
    2.6901e-06, 2.5853e-06, 2.5167e-06, 2.4749e-06, 2.4425e-06, 2.4462e-06, 
    2.4654e-06, 2.4969e-06, 2.5456e-06, 2.6029e-06, 2.6919e-06, 2.7545e-06, 
    2.7946e-06, 2.8242e-06, 2.8406e-06, 2.8443e-06, 2.8455e-06, 2.8575e-06, 
    2.9031e-06, 2.9781e-06, 3.0894e-06, 3.2204e-06, 3.3812e-06, 3.5576e-06, 
    3.5734e-06, 3.5697e-06, 3.6737e-06, 3.9326e-06, 3.9449e-06, 3.8885e-06, 
    3.9707e-06, 4.0048e-06, 4.0022e-06, 3.8396e-06, 2.6041e-06,
  0.011688, 0.011369, 0.011235, 0.011154, 0.011095, 0.011044, 0.010987, 
    0.010875, 0.010744, 0.010569, 0.010303, 0.010206, 0.010103, 0.0097492, 
    0.0089967, 0.0037976, 0.0010022, 0.0010435, 0.0013313, 0.0013471, 
    0.001094, 0.00082967, 0.00082622, 0.0010802, 0.0012854, 0.00028056, 
    0.00010323, 5.3134e-05, 0.00014431, 0.00049478, 0.00082306, 0.00068282, 
    0.00041795, 0.00026033, 0.00025169, 0.00018238, 0.00011712, 8.3828e-05, 
    6.6138e-05, 4.4506e-05, 3.2036e-05, 2.3549e-05, 1.8674e-05, 1.5615e-05, 
    1.2865e-05, 1.0825e-05, 9.3066e-06, 1.0196e-05, 7.3535e-06, 5.3743e-06, 
    4.9255e-06, 4.1876e-06, 3.2745e-06, 3.2472e-06, 3.0798e-06, 2.8187e-06, 
    2.6897e-06, 2.5832e-06, 2.5119e-06, 2.4729e-06, 2.4422e-06, 2.4461e-06, 
    2.465e-06, 2.4961e-06, 2.5443e-06, 2.6015e-06, 2.6911e-06, 2.7538e-06, 
    2.7941e-06, 2.8244e-06, 2.8409e-06, 2.844e-06, 2.8453e-06, 2.858e-06, 
    2.9024e-06, 2.9784e-06, 3.0932e-06, 3.2205e-06, 3.381e-06, 3.549e-06, 
    3.5474e-06, 3.5492e-06, 3.6712e-06, 3.931e-06, 3.9447e-06, 3.8875e-06, 
    3.9725e-06, 4.0067e-06, 4.0047e-06, 3.823e-06, 2.5977e-06,
  0.011968, 0.011668, 0.011542, 0.011468, 0.011417, 0.011376, 0.011339, 
    0.011287, 0.011205, 0.011066, 0.010755, 0.010687, 0.010469, 0.0093545, 
    0.0088257, 0.0050029, 0.0010803, 0.0010975, 0.0013255, 0.001411, 
    0.0011446, 0.0009498, 0.0010241, 0.0014118, 0.0019556, 0.0003587, 
    8.6127e-05, 4.8273e-05, 0.00018328, 0.00060294, 0.00080765, 0.00067233, 
    0.00042828, 0.00027229, 0.00026148, 0.00018137, 0.00011042, 8.2018e-05, 
    6.4712e-05, 4.4666e-05, 3.2267e-05, 2.2983e-05, 1.7403e-05, 1.4509e-05, 
    1.2547e-05, 1.0887e-05, 9.445e-06, 9.3096e-06, 7.4418e-06, 5.4884e-06, 
    5.1366e-06, 4.2457e-06, 3.2431e-06, 3.2251e-06, 3.078e-06, 2.8165e-06, 
    2.6876e-06, 2.5813e-06, 2.5082e-06, 2.4705e-06, 2.4421e-06, 2.4458e-06, 
    2.4644e-06, 2.4951e-06, 2.5428e-06, 2.6004e-06, 2.6902e-06, 2.7536e-06, 
    2.794e-06, 2.8247e-06, 2.8412e-06, 2.8437e-06, 2.845e-06, 2.8584e-06, 
    2.9019e-06, 2.9787e-06, 3.096e-06, 3.2202e-06, 3.3824e-06, 3.5399e-06, 
    3.5214e-06, 3.5292e-06, 3.6701e-06, 3.9281e-06, 3.9437e-06, 3.8865e-06, 
    3.9743e-06, 4.0091e-06, 4.0078e-06, 3.8063e-06, 2.5912e-06,
  0.012156, 0.011863, 0.011739, 0.011665, 0.011618, 0.011581, 0.011553, 
    0.011525, 0.011453, 0.011369, 0.011066, 0.011164, 0.010885, 0.0092056, 
    0.0090105, 0.0062258, 0.0012278, 0.0012313, 0.0013239, 0.0014854, 
    0.0012232, 0.0011058, 0.0012329, 0.0018066, 0.0026903, 0.00046334, 
    6.899e-05, 4.586e-05, 0.0001974, 0.00068275, 0.00078404, 0.00065911, 
    0.00043889, 0.00028201, 0.00026788, 0.00017763, 0.00010365, 8.1468e-05, 
    6.3889e-05, 4.5118e-05, 3.2462e-05, 2.2443e-05, 1.6198e-05, 1.3595e-05, 
    1.2293e-05, 1.0863e-05, 9.7913e-06, 8.4763e-06, 7.4673e-06, 5.5729e-06, 
    5.3565e-06, 4.2925e-06, 3.2143e-06, 3.2097e-06, 3.0782e-06, 2.8151e-06, 
    2.6858e-06, 2.5787e-06, 2.5046e-06, 2.4685e-06, 2.4422e-06, 2.4454e-06, 
    2.4638e-06, 2.4939e-06, 2.5412e-06, 2.5993e-06, 2.6893e-06, 2.7535e-06, 
    2.794e-06, 2.825e-06, 2.8414e-06, 2.8434e-06, 2.8447e-06, 2.8587e-06, 
    2.9017e-06, 2.9793e-06, 3.0985e-06, 3.2195e-06, 3.3842e-06, 3.5304e-06, 
    3.494e-06, 3.5089e-06, 3.6688e-06, 3.9249e-06, 3.9425e-06, 3.8854e-06, 
    3.976e-06, 4.0115e-06, 4.0108e-06, 3.79e-06, 2.5846e-06,
  0.0123, 0.012005, 0.011879, 0.011804, 0.011754, 0.011718, 0.011686, 
    0.011643, 0.011533, 0.011396, 0.011118, 0.011349, 0.011, 0.0093365, 
    0.0091656, 0.0073202, 0.0017738, 0.0013596, 0.0013581, 0.0015894, 
    0.0013903, 0.0013113, 0.0015215, 0.0023618, 0.0032923, 0.00074444, 
    6.3836e-05, 8.6519e-05, 0.00027242, 0.00071138, 0.00074426, 0.00062004, 
    0.00043635, 0.0002894, 0.00026015, 0.00016966, 0.00010133, 8.2601e-05, 
    6.3773e-05, 4.6086e-05, 3.2438e-05, 2.2215e-05, 1.5483e-05, 1.3423e-05, 
    1.2378e-05, 1.0959e-05, 1.0144e-05, 8.4214e-06, 7.4121e-06, 5.5604e-06, 
    5.1125e-06, 4.3047e-06, 3.1926e-06, 3.1924e-06, 3.0741e-06, 2.8136e-06, 
    2.6825e-06, 2.575e-06, 2.4999e-06, 2.465e-06, 2.4421e-06, 2.4448e-06, 
    2.4628e-06, 2.4926e-06, 2.5395e-06, 2.5991e-06, 2.6888e-06, 2.7532e-06, 
    2.794e-06, 2.8251e-06, 2.8415e-06, 2.8432e-06, 2.8446e-06, 2.859e-06, 
    2.9021e-06, 2.981e-06, 3.0995e-06, 3.2172e-06, 3.386e-06, 3.5176e-06, 
    3.466e-06, 3.4926e-06, 3.6625e-06, 3.9204e-06, 3.9411e-06, 3.8849e-06, 
    3.9774e-06, 4.0142e-06, 4.013e-06, 3.779e-06, 2.5766e-06,
  0.0124, 0.012104, 0.011979, 0.011904, 0.011854, 0.011819, 0.011789, 
    0.01175, 0.011652, 0.011507, 0.01118, 0.011438, 0.01108, 0.009698, 
    0.0090983, 0.0077231, 0.0023566, 0.001476, 0.0014032, 0.0017104, 
    0.001583, 0.0015223, 0.0018307, 0.0029439, 0.0038514, 0.0011425, 
    7.0825e-05, 0.0001315, 0.00042205, 0.00072199, 0.00070307, 0.00057984, 
    0.00043311, 0.00029622, 0.00024819, 0.00016113, 0.00010116, 8.4197e-05, 
    6.3774e-05, 4.7112e-05, 3.2305e-05, 2.1962e-05, 1.5016e-05, 1.3449e-05, 
    1.253e-05, 1.1178e-05, 1.0274e-05, 8.7249e-06, 7.3786e-06, 5.4751e-06, 
    4.8249e-06, 4.3086e-06, 3.1787e-06, 3.1792e-06, 3.069e-06, 2.8123e-06, 
    2.6803e-06, 2.5717e-06, 2.4953e-06, 2.4618e-06, 2.442e-06, 2.4444e-06, 
    2.462e-06, 2.4912e-06, 2.5381e-06, 2.5991e-06, 2.6882e-06, 2.7528e-06, 
    2.7938e-06, 2.8252e-06, 2.8416e-06, 2.8431e-06, 2.8444e-06, 2.8592e-06, 
    2.9025e-06, 2.9827e-06, 3.0997e-06, 3.2147e-06, 3.3876e-06, 3.5035e-06, 
    3.4413e-06, 3.4799e-06, 3.654e-06, 3.9151e-06, 3.9396e-06, 3.8843e-06, 
    3.9785e-06, 4.0165e-06, 4.0149e-06, 3.7713e-06, 2.5682e-06,
  0.01254, 0.012252, 0.012129, 0.012056, 0.012007, 0.011972, 0.011944, 
    0.011912, 0.011819, 0.011627, 0.011282, 0.011455, 0.011165, 0.010077, 
    0.0091711, 0.0075037, 0.0028142, 0.0016516, 0.0014704, 0.0018144, 
    0.0017498, 0.0017047, 0.0020584, 0.0033743, 0.0042751, 0.0017229, 
    0.00015236, 0.00021064, 0.00062545, 0.0007108, 0.00066556, 0.00054535, 
    0.00042822, 0.00030277, 0.00023448, 0.00015172, 0.00010308, 8.4822e-05, 
    6.4006e-05, 4.7784e-05, 3.2256e-05, 2.1612e-05, 1.4828e-05, 1.362e-05, 
    1.271e-05, 1.149e-05, 1.0207e-05, 9.2662e-06, 7.4992e-06, 5.3898e-06, 
    4.6352e-06, 4.2817e-06, 3.1745e-06, 3.1653e-06, 3.0615e-06, 2.8136e-06, 
    2.6795e-06, 2.5688e-06, 2.4906e-06, 2.4591e-06, 2.442e-06, 2.4442e-06, 
    2.4615e-06, 2.4899e-06, 2.537e-06, 2.5991e-06, 2.6875e-06, 2.7523e-06, 
    2.7937e-06, 2.8254e-06, 2.8416e-06, 2.843e-06, 2.8442e-06, 2.8594e-06, 
    2.9027e-06, 2.984e-06, 3.0994e-06, 3.2128e-06, 3.3887e-06, 3.4873e-06, 
    3.4221e-06, 3.4736e-06, 3.6443e-06, 3.9096e-06, 3.938e-06, 3.8835e-06, 
    3.9793e-06, 4.0181e-06, 4.0168e-06, 3.7677e-06, 2.5597e-06,
  0.012696, 0.012418, 0.0123, 0.012229, 0.01218, 0.012144, 0.012116, 
    0.012078, 0.011954, 0.011678, 0.011333, 0.011434, 0.011214, 0.010162, 
    0.0094889, 0.0073368, 0.0032488, 0.001877, 0.00152, 0.0018765, 0.0018602, 
    0.0018484, 0.0021714, 0.0036401, 0.0045685, 0.0024368, 0.00033215, 
    0.00033244, 0.00078716, 0.00068973, 0.00062959, 0.00051602, 0.00041967, 
    0.00030931, 0.00022129, 0.00014257, 0.00010638, 8.4721e-05, 6.4617e-05, 
    4.7847e-05, 3.221e-05, 2.1082e-05, 1.4888e-05, 1.3945e-05, 1.2939e-05, 
    1.1829e-05, 1.0159e-05, 9.7417e-06, 7.6656e-06, 5.4119e-06, 4.5377e-06, 
    4.182e-06, 3.1842e-06, 3.1543e-06, 3.0523e-06, 2.8139e-06, 2.6783e-06, 
    2.566e-06, 2.4858e-06, 2.4568e-06, 2.442e-06, 2.4443e-06, 2.4615e-06, 
    2.489e-06, 2.5363e-06, 2.5993e-06, 2.6864e-06, 2.7515e-06, 2.7935e-06, 
    2.8257e-06, 2.8416e-06, 2.843e-06, 2.844e-06, 2.8596e-06, 2.9025e-06, 
    2.9846e-06, 3.0988e-06, 3.2124e-06, 3.3893e-06, 3.4692e-06, 3.4092e-06, 
    3.4731e-06, 3.6333e-06, 3.9041e-06, 3.9362e-06, 3.883e-06, 3.9799e-06, 
    4.0191e-06, 4.0184e-06, 3.7669e-06, 2.552e-06,
  0.012943, 0.012679, 0.012567, 0.012499, 0.012452, 0.012417, 0.01239, 
    0.012351, 0.012221, 0.011877, 0.011691, 0.011598, 0.011112, 0.010082, 
    0.0096713, 0.0075222, 0.0036725, 0.0021989, 0.0015298, 0.0018525, 
    0.0018961, 0.0019679, 0.0022022, 0.0037149, 0.0046551, 0.0030226, 
    0.00071043, 0.00056636, 0.00082449, 0.00067515, 0.00059401, 0.00049498, 
    0.00041489, 0.00030931, 0.00020838, 0.00013297, 0.00010855, 8.4864e-05, 
    6.5852e-05, 4.7212e-05, 3.225e-05, 2.0404e-05, 1.5158e-05, 1.4387e-05, 
    1.3194e-05, 1.2036e-05, 1.0317e-05, 9.6262e-06, 7.8557e-06, 5.608e-06, 
    4.5565e-06, 3.9007e-06, 3.1974e-06, 3.1535e-06, 3.0325e-06, 2.8162e-06, 
    2.6776e-06, 2.5644e-06, 2.4823e-06, 2.4546e-06, 2.4418e-06, 2.4445e-06, 
    2.462e-06, 2.4894e-06, 2.5364e-06, 2.5995e-06, 2.6849e-06, 2.7502e-06, 
    2.7931e-06, 2.8258e-06, 2.8416e-06, 2.8429e-06, 2.844e-06, 2.8599e-06, 
    2.9017e-06, 2.9847e-06, 3.0983e-06, 3.2135e-06, 3.3894e-06, 3.4496e-06, 
    3.4002e-06, 3.4765e-06, 3.6216e-06, 3.8985e-06, 3.9346e-06, 3.8832e-06, 
    3.9806e-06, 4.0194e-06, 4.0194e-06, 3.7658e-06, 2.5467e-06,
  0.013209, 0.012959, 0.012852, 0.012787, 0.012741, 0.012708, 0.012678, 
    0.012625, 0.012501, 0.01204, 0.012067, 0.011761, 0.011017, 0.0099407, 
    0.0095998, 0.0078567, 0.0041381, 0.0026073, 0.0015344, 0.0017784, 
    0.0019058, 0.0020825, 0.0022238, 0.0036772, 0.0046176, 0.0034386, 
    0.0012081, 0.0008247, 0.00080948, 0.00066262, 0.00056317, 0.00048659, 
    0.00041501, 0.00030229, 0.00019577, 0.00012348, 0.00011028, 8.595e-05, 
    6.7e-05, 4.6372e-05, 3.2334e-05, 1.9637e-05, 1.5435e-05, 1.475e-05, 
    1.3362e-05, 1.213e-05, 1.0471e-05, 9.2264e-06, 8.0364e-06, 5.8538e-06, 
    4.6138e-06, 3.6652e-06, 3.1979e-06, 3.1602e-06, 3.0114e-06, 2.8173e-06, 
    2.6771e-06, 2.5638e-06, 2.4794e-06, 2.4525e-06, 2.4416e-06, 2.4447e-06, 
    2.4627e-06, 2.4902e-06, 2.5368e-06, 2.5995e-06, 2.683e-06, 2.7488e-06, 
    2.7928e-06, 2.8261e-06, 2.8416e-06, 2.8428e-06, 2.8442e-06, 2.8601e-06, 
    2.9004e-06, 2.985e-06, 3.0983e-06, 3.2159e-06, 3.3895e-06, 3.4304e-06, 
    3.39e-06, 3.4778e-06, 3.6103e-06, 3.8936e-06, 3.9327e-06, 3.8834e-06, 
    3.9813e-06, 4.0196e-06, 4.0201e-06, 3.7631e-06, 2.5421e-06,
  0.013496, 0.013263, 0.01316, 0.013097, 0.013053, 0.01302, 0.012983, 
    0.012906, 0.012748, 0.012259, 0.012309, 0.011788, 0.011079, 0.0099966, 
    0.0096464, 0.0083027, 0.004731, 0.0030344, 0.0015423, 0.0017071, 
    0.0019178, 0.0021892, 0.0022539, 0.0035695, 0.0045015, 0.0037245, 
    0.0016884, 0.0010231, 0.00082553, 0.00065037, 0.00053711, 0.00048328, 
    0.00040872, 0.00028569, 0.00018215, 0.00011752, 0.00011257, 8.8202e-05, 
    6.6865e-05, 4.5721e-05, 3.2437e-05, 1.8822e-05, 1.5701e-05, 1.5024e-05, 
    1.3413e-05, 1.2131e-05, 1.053e-05, 8.8729e-06, 8.0659e-06, 6.0581e-06, 
    4.6851e-06, 3.5537e-06, 3.1891e-06, 3.1688e-06, 2.9906e-06, 2.8152e-06, 
    2.6765e-06, 2.5637e-06, 2.477e-06, 2.4507e-06, 2.4413e-06, 2.4448e-06, 
    2.4633e-06, 2.4913e-06, 2.5377e-06, 2.5994e-06, 2.6808e-06, 2.7473e-06, 
    2.7927e-06, 2.8266e-06, 2.8416e-06, 2.8426e-06, 2.8445e-06, 2.8602e-06, 
    2.8987e-06, 2.9854e-06, 3.0986e-06, 3.2187e-06, 3.3895e-06, 3.413e-06, 
    3.3792e-06, 3.4747e-06, 3.5988e-06, 3.8891e-06, 3.9306e-06, 3.8835e-06, 
    3.9822e-06, 4.0195e-06, 4.0205e-06, 3.7579e-06, 2.5382e-06,
  0.013789, 0.013577, 0.013479, 0.01342, 0.013378, 0.013346, 0.013295, 
    0.013203, 0.012909, 0.012725, 0.012548, 0.011761, 0.011224, 0.01032, 
    0.01, 0.00913, 0.0055914, 0.003547, 0.001652, 0.0016781, 0.0019318, 
    0.0022576, 0.00227, 0.0033569, 0.0042576, 0.0038325, 0.0020065, 
    0.0011295, 0.00089402, 0.00064285, 0.00051674, 0.00048218, 0.00039485, 
    0.00025221, 0.00016364, 0.00011815, 0.00011509, 9.0181e-05, 6.496e-05, 
    4.5536e-05, 3.2413e-05, 1.8206e-05, 1.5961e-05, 1.5144e-05, 1.3209e-05, 
    1.1968e-05, 1.0368e-05, 8.6392e-06, 7.8122e-06, 6.1592e-06, 4.7524e-06, 
    3.497e-06, 3.1843e-06, 3.175e-06, 2.971e-06, 2.8149e-06, 2.6738e-06, 
    2.5638e-06, 2.476e-06, 2.4491e-06, 2.4408e-06, 2.4447e-06, 2.464e-06, 
    2.4927e-06, 2.5386e-06, 2.5992e-06, 2.6785e-06, 2.746e-06, 2.793e-06, 
    2.8271e-06, 2.8416e-06, 2.8425e-06, 2.8451e-06, 2.8605e-06, 2.8967e-06, 
    2.9857e-06, 3.0982e-06, 3.2215e-06, 3.3895e-06, 3.3997e-06, 3.3694e-06, 
    3.4652e-06, 3.5889e-06, 3.8851e-06, 3.9285e-06, 3.8833e-06, 3.9828e-06, 
    4.0186e-06, 4.0199e-06, 3.7477e-06, 2.5339e-06,
  0.014031, 0.013836, 0.013743, 0.013687, 0.013646, 0.013608, 0.013538, 
    0.013424, 0.013039, 0.013106, 0.012704, 0.011818, 0.011379, 0.010542, 
    0.01023, 0.0096929, 0.0063452, 0.0041792, 0.0019207, 0.0016861, 
    0.0019438, 0.0023056, 0.0022672, 0.003143, 0.0040271, 0.0038722, 
    0.0022266, 0.0012191, 0.0009529, 0.00063701, 0.00050055, 0.00047857, 
    0.00037617, 0.00021692, 0.00014373, 0.00012096, 0.00011701, 9e-05, 
    6.2501e-05, 4.5385e-05, 3.1827e-05, 1.7836e-05, 1.6233e-05, 1.5222e-05, 
    1.2865e-05, 1.1634e-05, 1.0142e-05, 8.3807e-06, 7.5109e-06, 6.1909e-06, 
    4.8282e-06, 3.438e-06, 3.193e-06, 3.1787e-06, 2.9553e-06, 2.8117e-06, 
    2.6704e-06, 2.5637e-06, 2.4755e-06, 2.4477e-06, 2.4403e-06, 2.4444e-06, 
    2.4645e-06, 2.4941e-06, 2.5396e-06, 2.599e-06, 2.6761e-06, 2.7448e-06, 
    2.7936e-06, 2.8275e-06, 2.8417e-06, 2.8425e-06, 2.846e-06, 2.8608e-06, 
    2.8949e-06, 2.9855e-06, 3.0965e-06, 3.2241e-06, 3.3895e-06, 3.3892e-06, 
    3.3619e-06, 3.4523e-06, 3.58e-06, 3.8808e-06, 3.9266e-06, 3.8827e-06, 
    3.9832e-06, 4.0168e-06, 4.0183e-06, 3.7348e-06, 2.5279e-06,
  0.014247, 0.014066, 0.013978, 0.013922, 0.013878, 0.013831, 0.013731, 
    0.013523, 0.013193, 0.013202, 0.012754, 0.01192, 0.011426, 0.010622, 
    0.010231, 0.0098195, 0.0070163, 0.0048037, 0.0023757, 0.0017609, 
    0.0019612, 0.0023295, 0.0022474, 0.00298, 0.0038251, 0.0037811, 
    0.0023278, 0.0013117, 0.00097278, 0.00063577, 0.0004972, 0.00047705, 
    0.00035531, 0.00018674, 0.00012673, 0.00012339, 0.00011664, 8.655e-05, 
    6.0029e-05, 4.5441e-05, 3.09e-05, 1.7723e-05, 1.6546e-05, 1.5418e-05, 
    1.2553e-05, 1.1124e-05, 9.937e-06, 8.1527e-06, 7.1801e-06, 6.1021e-06, 
    4.895e-06, 3.3641e-06, 3.2007e-06, 3.1703e-06, 2.9435e-06, 2.8071e-06, 
    2.6671e-06, 2.5635e-06, 2.475e-06, 2.4465e-06, 2.4398e-06, 2.4441e-06, 
    2.4647e-06, 2.4952e-06, 2.5407e-06, 2.5988e-06, 2.6738e-06, 2.7438e-06, 
    2.794e-06, 2.8279e-06, 2.8418e-06, 2.8426e-06, 2.8472e-06, 2.8614e-06, 
    2.8936e-06, 2.9849e-06, 3.0934e-06, 3.2256e-06, 3.3891e-06, 3.382e-06, 
    3.3566e-06, 3.4367e-06, 3.5726e-06, 3.8761e-06, 3.9242e-06, 3.8812e-06, 
    3.9836e-06, 4.0146e-06, 4.016e-06, 3.7206e-06, 2.5208e-06,
  0.014475, 0.014312, 0.014228, 0.014171, 0.014123, 0.014072, 0.013948, 
    0.013619, 0.013357, 0.013257, 0.012839, 0.011987, 0.011409, 0.010678, 
    0.010231, 0.0099932, 0.0079119, 0.0054415, 0.0028505, 0.0018446, 
    0.0019819, 0.0023433, 0.0022215, 0.0028555, 0.0036583, 0.003683, 
    0.002403, 0.0014029, 0.00099288, 0.00064113, 0.00049651, 0.00047453, 
    0.00033723, 0.00016389, 0.00011546, 0.00012413, 0.00011541, 8.2493e-05, 
    5.8028e-05, 4.5293e-05, 2.9648e-05, 1.7679e-05, 1.6873e-05, 1.5669e-05, 
    1.2293e-05, 1.051e-05, 9.7227e-06, 7.9441e-06, 6.8924e-06, 6.0046e-06, 
    4.9409e-06, 3.2906e-06, 3.2256e-06, 3.16e-06, 2.9369e-06, 2.8006e-06, 
    2.662e-06, 2.5628e-06, 2.4738e-06, 2.4455e-06, 2.4393e-06, 2.4437e-06, 
    2.4647e-06, 2.4962e-06, 2.5419e-06, 2.5986e-06, 2.6714e-06, 2.7429e-06, 
    2.7945e-06, 2.8286e-06, 2.8418e-06, 2.8427e-06, 2.8486e-06, 2.8622e-06, 
    2.8926e-06, 2.9839e-06, 3.0894e-06, 3.2274e-06, 3.3886e-06, 3.3761e-06, 
    3.3526e-06, 3.4205e-06, 3.5658e-06, 3.8714e-06, 3.9213e-06, 3.8793e-06, 
    3.984e-06, 4.0122e-06, 4.0135e-06, 3.707e-06, 2.5123e-06,
  0.014479, 0.014314, 0.014233, 0.014179, 0.014131, 0.014064, 0.013938, 
    0.013504, 0.013134, 0.012932, 0.012551, 0.011899, 0.011353, 0.010753, 
    0.010229, 0.0098666, 0.0086731, 0.0060086, 0.0032269, 0.0020284, 
    0.0020443, 0.0023347, 0.0022062, 0.002828, 0.0035613, 0.0036174, 
    0.0024871, 0.0014999, 0.0010026, 0.00065457, 0.00050707, 0.00047345, 
    0.00032305, 0.00015733, 0.0001149, 0.00012025, 0.00011032, 7.8043e-05, 
    5.7649e-05, 4.4727e-05, 2.8054e-05, 1.7953e-05, 1.7391e-05, 1.631e-05, 
    1.2558e-05, 9.9806e-06, 9.3252e-06, 7.9552e-06, 6.7955e-06, 6.0038e-06, 
    4.8912e-06, 3.1998e-06, 3.2577e-06, 3.1501e-06, 2.9422e-06, 2.796e-06, 
    2.66e-06, 2.5618e-06, 2.474e-06, 2.4445e-06, 2.4389e-06, 2.4437e-06, 
    2.4649e-06, 2.4964e-06, 2.5427e-06, 2.5985e-06, 2.6694e-06, 2.742e-06, 
    2.7949e-06, 2.8292e-06, 2.8419e-06, 2.8432e-06, 2.8505e-06, 2.8638e-06, 
    2.8928e-06, 2.9815e-06, 3.0841e-06, 3.2279e-06, 3.3867e-06, 3.3727e-06, 
    3.3533e-06, 3.4095e-06, 3.5658e-06, 3.8631e-06, 3.9178e-06, 3.8768e-06, 
    3.9843e-06, 4.0106e-06, 4.0115e-06, 3.6937e-06, 2.5022e-06,
  0.014543, 0.014381, 0.0143, 0.014246, 0.014201, 0.014115, 0.013969, 
    0.013381, 0.012892, 0.012642, 0.012334, 0.011894, 0.011421, 0.010866, 
    0.010254, 0.0098514, 0.009449, 0.0067898, 0.0036314, 0.0023076, 0.002132, 
    0.0023222, 0.0022045, 0.0028196, 0.0034743, 0.0035382, 0.0025276, 
    0.0015761, 0.0010142, 0.00067118, 0.00051974, 0.00047489, 0.00031318, 
    0.00015255, 0.00011491, 0.00011667, 0.00010412, 7.4065e-05, 5.7379e-05, 
    4.3841e-05, 2.6453e-05, 1.8212e-05, 1.7982e-05, 1.7023e-05, 1.2926e-05, 
    9.586e-06, 8.9398e-06, 7.9294e-06, 6.7211e-06, 6.0117e-06, 4.8284e-06, 
    3.1187e-06, 3.291e-06, 3.1467e-06, 2.9506e-06, 2.7899e-06, 2.6578e-06, 
    2.5607e-06, 2.4738e-06, 2.4439e-06, 2.4386e-06, 2.4438e-06, 2.4651e-06, 
    2.4964e-06, 2.5435e-06, 2.5982e-06, 2.6676e-06, 2.7411e-06, 2.7953e-06, 
    2.8298e-06, 2.842e-06, 2.8437e-06, 2.8524e-06, 2.8656e-06, 2.8934e-06, 
    2.979e-06, 3.0792e-06, 3.2289e-06, 3.3843e-06, 3.3689e-06, 3.355e-06, 
    3.4007e-06, 3.5672e-06, 3.8538e-06, 3.914e-06, 3.8746e-06, 3.9845e-06, 
    4.0091e-06, 4.0095e-06, 3.6811e-06, 2.4921e-06,
  0.014588, 0.014433, 0.014353, 0.014298, 0.014255, 0.014185, 0.014068, 
    0.013397, 0.01291, 0.012683, 0.012354, 0.011932, 0.011468, 0.010905, 
    0.010235, 0.0099136, 0.0097137, 0.0074644, 0.0040027, 0.0026316, 
    0.0022383, 0.0022969, 0.0022234, 0.0028491, 0.0034727, 0.003476, 
    0.0025512, 0.0016272, 0.001039, 0.0006721, 0.00052713, 0.00046733, 
    0.00029764, 0.00015096, 0.00011625, 0.00011428, 9.6872e-05, 7.2319e-05, 
    5.7528e-05, 4.243e-05, 2.485e-05, 1.8427e-05, 1.8646e-05, 1.7828e-05, 
    1.3414e-05, 9.4371e-06, 8.6789e-06, 7.7581e-06, 6.7586e-06, 6.1517e-06, 
    4.7591e-06, 3.0501e-06, 3.3243e-06, 3.151e-06, 2.9594e-06, 2.78e-06, 
    2.6564e-06, 2.5594e-06, 2.4744e-06, 2.4435e-06, 2.4382e-06, 2.444e-06, 
    2.4652e-06, 2.4961e-06, 2.5437e-06, 2.5976e-06, 2.6662e-06, 2.7404e-06, 
    2.7954e-06, 2.8303e-06, 2.8422e-06, 2.8443e-06, 2.854e-06, 2.8673e-06, 
    2.8946e-06, 2.9767e-06, 3.0751e-06, 3.2292e-06, 3.3829e-06, 3.3647e-06, 
    3.3577e-06, 3.3948e-06, 3.5679e-06, 3.8416e-06, 3.91e-06, 3.8732e-06, 
    3.9845e-06, 4.0078e-06, 4.0075e-06, 3.6683e-06, 2.4818e-06,
  0.014594, 0.014448, 0.014373, 0.014322, 0.014281, 0.014237, 0.01417, 
    0.01348, 0.013032, 0.012809, 0.012459, 0.011996, 0.011529, 0.010962, 
    0.010233, 0.010014, 0.0099622, 0.0079903, 0.0043318, 0.0029135, 
    0.0023356, 0.0022615, 0.0022499, 0.0028815, 0.0034754, 0.0034287, 
    0.0025691, 0.0016734, 0.00106, 0.00067015, 0.00053431, 0.00046054, 
    0.00028178, 0.00014759, 0.00011599, 0.00011266, 9.0815e-05, 7.0967e-05, 
    5.7274e-05, 4.0795e-05, 2.3392e-05, 1.8644e-05, 1.9395e-05, 1.8675e-05, 
    1.3865e-05, 9.3718e-06, 8.5915e-06, 7.5988e-06, 6.76e-06, 6.267e-06, 
    4.6943e-06, 2.9906e-06, 3.3525e-06, 3.1617e-06, 2.9709e-06, 2.7709e-06, 
    2.6537e-06, 2.558e-06, 2.4749e-06, 2.4433e-06, 2.438e-06, 2.4442e-06, 
    2.4653e-06, 2.4958e-06, 2.5439e-06, 2.5966e-06, 2.665e-06, 2.7398e-06, 
    2.7954e-06, 2.831e-06, 2.8425e-06, 2.8448e-06, 2.8555e-06, 2.869e-06, 
    2.8958e-06, 2.9749e-06, 3.0716e-06, 3.2297e-06, 3.3812e-06, 3.3594e-06, 
    3.36e-06, 3.3899e-06, 3.5677e-06, 3.8279e-06, 3.9059e-06, 3.8723e-06, 
    3.9847e-06, 4.0067e-06, 4.0055e-06, 3.6573e-06, 2.4716e-06,
  0.014635, 0.014489, 0.014417, 0.014363, 0.01432, 0.014264, 0.014105, 
    0.01349, 0.013138, 0.012952, 0.012616, 0.012082, 0.011481, 0.010857, 
    0.010217, 0.0099475, 0.0099533, 0.0080103, 0.004668, 0.0031752, 0.002404, 
    0.002234, 0.0022898, 0.0029283, 0.0034948, 0.0033697, 0.0025421, 
    0.0017093, 0.0010587, 0.00066767, 0.00053277, 0.00044216, 0.00026375, 
    0.00014577, 0.00011435, 0.00011376, 9.2456e-05, 7.0844e-05, 5.6043e-05, 
    3.8451e-05, 2.262e-05, 1.919e-05, 2.0317e-05, 1.9543e-05, 1.4342e-05, 
    9.524e-06, 8.6311e-06, 7.6406e-06, 6.7263e-06, 6.2637e-06, 4.6412e-06, 
    2.946e-06, 3.3308e-06, 3.1779e-06, 2.9715e-06, 2.7611e-06, 2.6506e-06, 
    2.5586e-06, 2.478e-06, 2.4426e-06, 2.4381e-06, 2.4449e-06, 2.4655e-06, 
    2.4953e-06, 2.5431e-06, 2.5953e-06, 2.6646e-06, 2.7389e-06, 2.7944e-06, 
    2.8314e-06, 2.843e-06, 2.8456e-06, 2.8563e-06, 2.8704e-06, 2.8968e-06, 
    2.974e-06, 3.0689e-06, 3.2299e-06, 3.3782e-06, 3.3533e-06, 3.359e-06, 
    3.388e-06, 3.567e-06, 3.812e-06, 3.9018e-06, 3.8713e-06, 3.9859e-06, 
    4.0073e-06, 4.0053e-06, 3.6539e-06, 2.4616e-06,
  0.014682, 0.014537, 0.014465, 0.014412, 0.014372, 0.014296, 0.014069, 
    0.013479, 0.013207, 0.013063, 0.012744, 0.012156, 0.011441, 0.010755, 
    0.010169, 0.009827, 0.0098559, 0.0078453, 0.0049572, 0.0034364, 
    0.0024876, 0.0022239, 0.0023309, 0.0029864, 0.0035106, 0.0033116, 
    0.0025255, 0.0017443, 0.001046, 0.00066354, 0.00052988, 0.00042421, 
    0.0002461, 0.00014465, 0.00011274, 0.00011519, 9.595e-05, 7.0893e-05, 
    5.4425e-05, 3.5852e-05, 2.1975e-05, 1.9741e-05, 2.1276e-05, 2.035e-05, 
    1.4764e-05, 9.687e-06, 8.6232e-06, 7.6908e-06, 6.6749e-06, 6.202e-06, 
    4.5979e-06, 2.9095e-06, 3.2614e-06, 3.1941e-06, 2.9731e-06, 2.7497e-06, 
    2.6469e-06, 2.5594e-06, 2.481e-06, 2.4422e-06, 2.4382e-06, 2.4455e-06, 
    2.4657e-06, 2.495e-06, 2.5423e-06, 2.5937e-06, 2.6643e-06, 2.7382e-06, 
    2.7935e-06, 2.8319e-06, 2.8435e-06, 2.8463e-06, 2.857e-06, 2.8716e-06, 
    2.8976e-06, 2.9733e-06, 3.0662e-06, 3.2304e-06, 3.3751e-06, 3.3473e-06, 
    3.3555e-06, 3.3862e-06, 3.5645e-06, 3.7961e-06, 3.8974e-06, 3.8703e-06, 
    3.9876e-06, 4.0093e-06, 4.0066e-06, 3.6528e-06, 2.4515e-06,
  0.014713, 0.014573, 0.0145, 0.014452, 0.014415, 0.014319, 0.014023, 
    0.013404, 0.013201, 0.013061, 0.012757, 0.012155, 0.011401, 0.010684, 
    0.010084, 0.0097046, 0.009693, 0.0075696, 0.0051445, 0.0036706, 
    0.0025921, 0.0022432, 0.0023607, 0.0030292, 0.0034986, 0.0032655, 
    0.0025396, 0.0017606, 0.0010251, 0.00066341, 0.00052564, 0.00040703, 
    0.0002294, 0.0001437, 0.00011336, 0.00011738, 9.9411e-05, 7.0616e-05, 
    5.1797e-05, 3.2893e-05, 2.1469e-05, 2.0299e-05, 2.2266e-05, 2.1095e-05, 
    1.52e-05, 9.8563e-06, 8.5481e-06, 7.7278e-06, 6.6015e-06, 5.9975e-06, 
    4.5725e-06, 2.8813e-06, 3.1698e-06, 3.208e-06, 2.9687e-06, 2.7385e-06, 
    2.6419e-06, 2.5603e-06, 2.4838e-06, 2.4423e-06, 2.4381e-06, 2.4461e-06, 
    2.4656e-06, 2.4946e-06, 2.5411e-06, 2.5919e-06, 2.6644e-06, 2.738e-06, 
    2.7928e-06, 2.8323e-06, 2.8441e-06, 2.8469e-06, 2.8577e-06, 2.8726e-06, 
    2.898e-06, 2.9723e-06, 3.0636e-06, 3.2315e-06, 3.372e-06, 3.3419e-06, 
    3.3477e-06, 3.3848e-06, 3.5599e-06, 3.7833e-06, 3.8934e-06, 3.8692e-06, 
    3.9898e-06, 4.0131e-06, 4.01e-06, 3.6537e-06, 2.4425e-06,
  0.014745, 0.014609, 0.014539, 0.01449, 0.014441, 0.014326, 0.013979, 
    0.013366, 0.013162, 0.012996, 0.012699, 0.012096, 0.011333, 0.010603, 
    0.010005, 0.0096034, 0.0094688, 0.007418, 0.0052026, 0.0038206, 
    0.0026743, 0.0022727, 0.0023889, 0.0030671, 0.0034798, 0.0032419, 
    0.0025803, 0.0017807, 0.0010117, 0.00066696, 0.00052237, 0.00039084, 
    0.00021273, 0.00014301, 0.00011568, 0.0001195, 0.00010033, 6.9697e-05, 
    4.8478e-05, 3.0065e-05, 2.1296e-05, 2.1086e-05, 2.3319e-05, 2.1706e-05, 
    1.5644e-05, 1.0009e-05, 8.3701e-06, 7.7201e-06, 6.4921e-06, 5.6743e-06, 
    4.5659e-06, 2.8592e-06, 3.0567e-06, 3.2168e-06, 2.9631e-06, 2.73e-06, 
    2.6369e-06, 2.5611e-06, 2.4863e-06, 2.4423e-06, 2.4382e-06, 2.4467e-06, 
    2.4655e-06, 2.4944e-06, 2.5398e-06, 2.5903e-06, 2.6646e-06, 2.7374e-06, 
    2.7919e-06, 2.8328e-06, 2.8447e-06, 2.8472e-06, 2.8584e-06, 2.8731e-06, 
    2.8981e-06, 2.9708e-06, 3.0614e-06, 3.2332e-06, 3.3694e-06, 3.3376e-06, 
    3.3373e-06, 3.3841e-06, 3.5525e-06, 3.7723e-06, 3.8889e-06, 3.8689e-06, 
    3.9925e-06, 4.0195e-06, 4.0162e-06, 3.6524e-06, 2.4374e-06,
  0.014764, 0.014632, 0.014564, 0.014507, 0.014426, 0.014277, 0.013943, 
    0.013332, 0.013061, 0.012856, 0.012539, 0.011956, 0.011214, 0.010507, 
    0.0099455, 0.0094434, 0.0091868, 0.007197, 0.0052642, 0.0039213, 
    0.0027043, 0.0022844, 0.0024192, 0.0031111, 0.003481, 0.0032239, 
    0.0026122, 0.001813, 0.0010148, 0.00067064, 0.00052129, 0.00037491, 
    0.00019867, 0.00014234, 0.0001186, 0.00012051, 9.7978e-05, 6.7191e-05, 
    4.4528e-05, 2.7831e-05, 2.1432e-05, 2.2318e-05, 2.4471e-05, 2.2295e-05, 
    1.6224e-05, 1.0278e-05, 8.1057e-06, 7.5607e-06, 6.3905e-06, 5.3466e-06, 
    4.5508e-06, 2.8463e-06, 3.0063e-06, 3.2204e-06, 2.9594e-06, 2.7214e-06, 
    2.6324e-06, 2.5613e-06, 2.4886e-06, 2.4422e-06, 2.4383e-06, 2.4472e-06, 
    2.4653e-06, 2.4942e-06, 2.5383e-06, 2.5891e-06, 2.6649e-06, 2.7364e-06, 
    2.7907e-06, 2.8331e-06, 2.8452e-06, 2.8475e-06, 2.8591e-06, 2.873e-06, 
    2.8979e-06, 2.9687e-06, 3.0605e-06, 3.2358e-06, 3.3668e-06, 3.3346e-06, 
    3.3269e-06, 3.3838e-06, 3.5413e-06, 3.7637e-06, 3.8842e-06, 3.8694e-06, 
    3.9946e-06, 4.0269e-06, 4.0235e-06, 3.6453e-06, 2.4372e-06,
  0.014765, 0.014635, 0.01457, 0.014509, 0.01439, 0.01419, 0.013899, 
    0.013323, 0.012975, 0.012722, 0.012389, 0.011824, 0.011102, 0.010428, 
    0.0099221, 0.0093403, 0.0089994, 0.0069125, 0.0053555, 0.0040363, 
    0.0027209, 0.0022817, 0.0024422, 0.0031616, 0.0034982, 0.003184, 
    0.0026172, 0.00185, 0.0010293, 0.00067525, 0.00052412, 0.00035848, 
    0.00018679, 0.00014136, 0.00012123, 0.00012087, 9.4281e-05, 6.3357e-05, 
    4.0041e-05, 2.5817e-05, 2.1578e-05, 2.375e-05, 2.5751e-05, 2.3061e-05, 
    1.6923e-05, 1.0701e-05, 7.8584e-06, 7.2621e-06, 6.341e-06, 5.1516e-06, 
    4.4705e-06, 2.8414e-06, 3.0428e-06, 3.2217e-06, 2.9544e-06, 2.711e-06, 
    2.628e-06, 2.5606e-06, 2.4907e-06, 2.4425e-06, 2.4385e-06, 2.4475e-06, 
    2.465e-06, 2.4939e-06, 2.5367e-06, 2.5882e-06, 2.6652e-06, 2.7353e-06, 
    2.7898e-06, 2.8334e-06, 2.8458e-06, 2.8479e-06, 2.8599e-06, 2.8729e-06, 
    2.8979e-06, 2.9664e-06, 3.0608e-06, 3.239e-06, 3.3633e-06, 3.3317e-06, 
    3.3173e-06, 3.3827e-06, 3.5282e-06, 3.7573e-06, 3.8799e-06, 3.8696e-06, 
    3.9961e-06, 4.0331e-06, 4.0298e-06, 3.6352e-06, 2.4387e-06 ;

 shum_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;

 meteo_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07 ;
}
