netcdf ropp_test_5o {
dimensions:
	dim_unlim = UNLIMITED ; // (2 currently)
	dim_char04 = 5 ;
	dim_char20 = 21 ;
	dim_char40 = 41 ;
	dim_char64 = 65 ;
	xyz = 3 ;
	dim_lev1b = 2319 ;
	dim_lev2a = 817 ;
variables:
	char occ_id(dim_unlim, dim_char40) ;
		occ_id:long_name = "Occultation ID" ;
	char gns_id(dim_unlim, dim_char04) ;
		gns_id:long_name = "GNSS satellite ID" ;
	char leo_id(dim_unlim, dim_char04) ;
		leo_id:long_name = "LEO satellite ID" ;
	char stn_id(dim_unlim, dim_char04) ;
		stn_id:long_name = "Ground station ID" ;
	double start_time(dim_unlim) ;
		start_time:long_name = "Starting time for the occultation" ;
		start_time:units = "seconds since 2000-01-01 00:00:00" ;
	int year(dim_unlim) ;
		year:long_name = "Year" ;
		year:units = "years" ;
		year:valid_range = 1995, 2099 ;
	int month(dim_unlim) ;
		month:long_name = "Month" ;
		month:units = "months" ;
		month:valid_range = 1, 12 ;
	int day(dim_unlim) ;
		day:long_name = "Day" ;
		day:units = "days" ;
		day:valid_range = 1, 31 ;
	int hour(dim_unlim) ;
		hour:long_name = "Hour" ;
		hour:units = "hours" ;
		hour:valid_range = 0, 23 ;
	int minute(dim_unlim) ;
		minute:long_name = "Minute" ;
		minute:units = "minutes" ;
		minute:valid_range = 0, 59 ;
	int second(dim_unlim) ;
		second:long_name = "Second" ;
		second:units = "seconds" ;
		second:valid_range = 0, 59 ;
	int msec(dim_unlim) ;
		msec:long_name = "Millisecond" ;
		msec:units = "milliseconds" ;
		msec:valid_range = 0, 999 ;
	int pcd(dim_unlim) ;
		pcd:long_name = "Product Confidence Data" ;
		pcd:units = "bits" ;
		pcd:valid_range = 0, 32767 ;
	float overall_qual(dim_unlim) ;
		overall_qual:long_name = "Overall quality" ;
		overall_qual:units = "percent" ;
		overall_qual:valid_range = 0., 100. ;
	double time(dim_unlim) ;
		time:long_name = "Reference time for the occultation" ;
		time:units = "seconds since 2000-01-01 00:00:00" ;
	float time_offset(dim_unlim) ;
		time_offset:long_name = "Time offset for georeferencing (since start of occ.)" ;
		time_offset:units = "seconds" ;
		time_offset:valid_range = 0., 240. ;
	float lat(dim_unlim) ;
		lat:long_name = "Reference latitude for the occultation" ;
		lat:units = "degrees_north" ;
		lat:valid_range = -90., 90. ;
	float lon(dim_unlim) ;
		lon:long_name = "Reference longitude for the occultation" ;
		lon:units = "degrees_east" ;
		lon:valid_range = -180., 180. ;
	float undulation(dim_unlim) ;
		undulation:long_name = "Geoid undulation for the reference coordinate" ;
		undulation:units = "metres" ;
		undulation:valid_range = -150., 150. ;
	double roc(dim_unlim) ;
		roc:long_name = "Radius of curvature for the reference coordinate" ;
		roc:units = "metres" ;
		roc:valid_range = 6.2e+06, 6.6e+06 ;
	float r_coc(dim_unlim, xyz) ;
		r_coc:long_name = "Centre of curvature for the reference coordinate" ;
		r_coc:units = "metres" ;
		r_coc:valid_range = -50000., 50000. ;
		r_coc:reference_frame = "ECF" ;
	float azimuth(dim_unlim) ;
		azimuth:long_name = "GNSS->LEO line of sight angle (from True North) for the reference coordinate" ;
		azimuth:units = "degrees_T" ;
		azimuth:valid_range = 0., 359.9 ;
	float lat_tp(dim_unlim, dim_lev1b) ;
		lat_tp:long_name = "Latitudes for tangent points" ;
		lat_tp:units = "degrees_north" ;
		lat_tp:valid_range = -90., 90. ;
	float lon_tp(dim_unlim, dim_lev1b) ;
		lon_tp:long_name = "Longitudes for tangent points" ;
		lon_tp:units = "degrees_east" ;
		lon_tp:valid_range = -180., 180. ;
	float azimuth_tp(dim_unlim, dim_lev1b) ;
		azimuth_tp:long_name = "GNSS->LEO line of sight angles (from True North) for tangent points" ;
		azimuth_tp:units = "degrees" ;
		azimuth_tp:valid_range = 0., 359.9 ;
	double impact_L1(dim_unlim, dim_lev1b) ;
		impact_L1:long_name = "Impact parameter (L1)" ;
		impact_L1:units = "metres" ;
		impact_L1:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_L2(dim_unlim, dim_lev1b) ;
		impact_L2:long_name = "Impact parameter (L2)" ;
		impact_L2:units = "metres" ;
		impact_L2:valid_range = 6.2e+06, 6.6e+06 ;
	double impact(dim_unlim, dim_lev1b) ;
		impact:long_name = "Impact parameter (generic)" ;
		impact:units = "metres" ;
		impact:valid_range = 6.2e+06, 6.6e+06 ;
	double impact_opt(dim_unlim, dim_lev1b) ;
		impact_opt:long_name = "Impact parameter (optimised)" ;
		impact_opt:units = "metres" ;
		impact_opt:valid_range = 6.2e+06, 6.6e+06 ;
	double bangle_L1(dim_unlim, dim_lev1b) ;
		bangle_L1:long_name = "Bending angle (L1)" ;
		bangle_L1:units = "radians" ;
		bangle_L1:valid_range = -0.001, 0.1 ;
	double bangle_L2(dim_unlim, dim_lev1b) ;
		bangle_L2:long_name = "Bending angle (L2)" ;
		bangle_L2:units = "radians" ;
		bangle_L2:valid_range = -0.001, 0.1 ;
	double bangle(dim_unlim, dim_lev1b) ;
		bangle:long_name = "Bending angle (generic)" ;
		bangle:units = "radians" ;
		bangle:valid_range = -0.001, 0.1 ;
	double bangle_opt(dim_unlim, dim_lev1b) ;
		bangle_opt:long_name = "Bending angle (optimised)" ;
		bangle_opt:units = "radians" ;
		bangle_opt:valid_range = -0.001, 0.1 ;
	double bangle_L1_sigma(dim_unlim, dim_lev1b) ;
		bangle_L1_sigma:long_name = "Estimated error (1-sigma) for bending angles (L1)" ;
		bangle_L1_sigma:units = "radians" ;
		bangle_L1_sigma:valid_range = 0., 0.01 ;
	double bangle_L2_sigma(dim_unlim, dim_lev1b) ;
		bangle_L2_sigma:long_name = "Estimated error (1-sigma) for bending angles (L2)" ;
		bangle_L2_sigma:units = "radians" ;
		bangle_L2_sigma:valid_range = 0., 0.01 ;
	double bangle_sigma(dim_unlim, dim_lev1b) ;
		bangle_sigma:long_name = "Estimated error (1-sigma) for bending angles (generic)" ;
		bangle_sigma:units = "radians" ;
		bangle_sigma:valid_range = 0., 0.01 ;
	double bangle_opt_sigma(dim_unlim, dim_lev1b) ;
		bangle_opt_sigma:long_name = "Estimated error (1-sigma) for bending angles (optimised)" ;
		bangle_opt_sigma:units = "radians" ;
		bangle_opt_sigma:valid_range = 0., 0.01 ;
	float bangle_L1_qual(dim_unlim, dim_lev1b) ;
		bangle_L1_qual:long_name = "Bending angle quality value (L1)" ;
		bangle_L1_qual:units = "percent" ;
		bangle_L1_qual:valid_range = 0., 100. ;
	float bangle_L2_qual(dim_unlim, dim_lev1b) ;
		bangle_L2_qual:long_name = "Bending angle quality value (L2)" ;
		bangle_L2_qual:units = "percent" ;
		bangle_L2_qual:valid_range = 0., 100. ;
	float bangle_qual(dim_unlim, dim_lev1b) ;
		bangle_qual:long_name = "Bending angle quality value (generic)" ;
		bangle_qual:units = "percent" ;
		bangle_qual:valid_range = 0., 100. ;
	float bangle_opt_qual(dim_unlim, dim_lev1b) ;
		bangle_opt_qual:long_name = "Bending angle quality value (optimised)" ;
		bangle_opt_qual:units = "percent" ;
		bangle_opt_qual:valid_range = 0., 100. ;
	float alt_refrac(dim_unlim, dim_lev2a) ;
		alt_refrac:long_name = "Geometric height above geoid for refractivity" ;
		alt_refrac:units = "metres" ;
		alt_refrac:valid_range = -1000., 1.e+05 ;
	float geop_refrac(dim_unlim, dim_lev2a) ;
		geop_refrac:long_name = "Geopotential height above geoid for refractivity" ;
		geop_refrac:units = "geopotential metres" ;
		geop_refrac:valid_range = -1000., 1.e+05 ;
	double refrac(dim_unlim, dim_lev2a) ;
		refrac:long_name = "Refractivity" ;
		refrac:units = "N-units" ;
		refrac:valid_range = 0., 500. ;
	double refrac_sigma(dim_unlim, dim_lev2a) ;
		refrac_sigma:long_name = "Estimated error (1-sigma) for refractivity" ;
		refrac_sigma:units = "N-units" ;
		refrac_sigma:valid_range = 0., 10. ;
	float refrac_qual(dim_unlim, dim_lev2a) ;
		refrac_qual:long_name = "Quality value for refractivity" ;
		refrac_qual:units = "percent" ;
		refrac_qual:valid_range = 0., 100. ;
	double dry_temp(dim_unlim, dim_lev2a) ;
		dry_temp:long_name = "Dry temperature" ;
		dry_temp:units = "kelvin" ;
		dry_temp:valid_range = 150., 350. ;
	double dry_temp_sigma(dim_unlim, dim_lev2a) ;
		dry_temp_sigma:long_name = "Estimated error (1-sigma) for dry temperature" ;
		dry_temp_sigma:units = "kelvin" ;
		dry_temp_sigma:valid_range = 0., 50. ;
	float dry_temp_qual(dim_unlim, dim_lev2a) ;
		dry_temp_qual:long_name = "Quality value for dry temperature" ;
		dry_temp_qual:units = "percent" ;
		dry_temp_qual:valid_range = 0., 100. ;

// global attributes:
		:title = "ROPP Radio Occultation data" ;
		:institution = "DMI GRAS SAF; Copyright 2009(C) EUMETSAT" ;
		:Conventions = "CF-1.0" ;
		:format_version = "ROPP I/O V1.1" ;
		:processing_centre = "DMI GRAS SAF; Copyright 2009(C) EUMETSAT" ;
		:processing_date = "2009-08-17 23:29:03.726" ;
		:pod_method = "UNDIFFERENCED Dynamical (SST)" ;
		:phase_method = "ND" ;
		:bangle_method = "GO" ;
		:refrac_method = "ABEL" ;
		:meteo_method = "1DV" ;
		:thin_method = "NONE (Thinning disabled) [v3.1]" ;
		:software_version = "UNKNOWN" ;
		:_FillValue = -9.9999e+07 ;
data:

 occ_id =
  "OC_20090817215807_META_G027_DMI_",
  "OC_20090817215807_META_G027_DMI_" ;

 gns_id =
  "G027",
  "G027" ;

 leo_id =
  "META",
  "META" ;

 stn_id =
  "NONE",
  "NONE" ;

 start_time = 3.0386e+08, 3.0386e+08 ;

 year = 2009, 2009 ;

 month = 8, 8 ;

 day = 17, 17 ;

 hour = 21, 21 ;

 minute = 58, 58 ;

 second = 7, 7 ;

 msec = 814, 814 ;

 pcd = 4, 4 ;

 overall_qual = -9.9999e+07, -9.9999e+07 ;

 time = 3.0386e+08, 3.0386e+08 ;

 time_offset = 5.7709, 5.7709 ;

 lat = 50.543, 50.543 ;

 lon = -3.89, -3.89 ;

 undulation = 52.499, 52.499 ;

 roc = 6.3745e+06, 6.3745e+06 ;

 r_coc =
  -3890.3, 9640.6, 20397,
  -3890.3, 9640.6, 20397 ;

 azimuth = -9.9999e+07, -9.9999e+07 ;

 lat_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 50.524, 50.524, 50.525, 50.525, 
    50.525, 50.526, 50.526, 50.527, 50.527, 50.527, 50.528, 50.528, 50.529, 
    50.529, 50.529, 50.53, 50.53, 50.531, 50.531, 50.531, 50.532, 50.532, 
    50.533, 50.533, 50.534, 50.534, 50.535, 50.535, 50.536, 50.536, 50.537, 
    50.537, 50.538, 50.538, 50.539, 50.54, 50.54, 50.541, 50.541, 50.542, 
    50.542, 50.543, 50.543, 50.544, 50.544, 50.544, 50.545, 50.545, 50.546, 
    50.546, 50.546, 50.547, 50.547, 50.547, 50.548, 50.548, 50.548, 50.549, 
    50.549, 50.549, 50.55, 50.55, 50.55, 50.551, 50.551, 50.551, 50.552, 
    50.552, 50.552, 50.553, 50.553, 50.553, 50.554, 50.554, 50.554, 50.555, 
    50.555, 50.555, 50.556, 50.556, 50.556, 50.557, 50.557, 50.557, 50.558, 
    50.558, 50.558, 50.559, 50.559, 50.56, 50.56, 50.56, 50.561, 50.561, 
    50.561, 50.562, 50.562, 50.563, 50.563, 50.563, 50.564, 50.564, 50.565, 
    50.565, 50.565, 50.566, 50.566, 50.567, 50.567, 50.567, 50.568, 50.568, 
    50.568, 50.569, 50.569, 50.57, 50.57, 50.57, 50.571, 50.571, 50.572, 
    50.572, 50.572, 50.573, 50.573, 50.573, 50.574, 50.574, 50.574, 50.575, 
    50.575, 50.575, 50.576, 50.576, 50.576, 50.577, 50.577, 50.577, 50.578, 
    50.578, 50.578, 50.579, 50.579, 50.579, 50.58, 50.58, 50.58, 50.58, 
    50.581, 50.581, 50.581, 50.581, 50.582, 50.582, 50.582, 50.583, 50.583, 
    50.583, 50.584, 50.584, 50.584, 50.584, 50.585, 50.585, 50.585, 50.586, 
    50.586, 50.586, 50.587, 50.587, 50.587, 50.588, 50.588, 50.588, 50.589, 
    50.589, 50.59, 50.59, 50.59, 50.591, 50.591, 50.591, 50.592, 50.592, 
    50.592, 50.593, 50.593, 50.593, 50.594, 50.594, 50.594, 50.595, 50.595, 
    50.595, 50.596, 50.596, 50.596, 50.597, 50.597, 50.597, 50.597, 50.598, 
    50.598, 50.598, 50.598, 50.599, 50.599, 50.599, 50.6, 50.6, 50.6, 50.6, 
    50.601, 50.601, 50.601, 50.602, 50.602, 50.602, 50.603, 50.603, 50.603, 
    50.604, 50.604, 50.604, 50.605, 50.605, 50.605, 50.606, 50.606, 50.606, 
    50.607, 50.607, 50.607, 50.607, 50.608, 50.608, 50.608, 50.608, 50.609, 
    50.609, 50.609, 50.61, 50.61, 50.61, 50.61, 50.61, 50.611, 50.611, 
    50.611, 50.612, 50.612, 50.612, 50.612, 50.613, 50.613, 50.613, 50.613, 
    50.614, 50.614, 50.614, 50.615, 50.615, 50.615, 50.615, 50.616, 50.616, 
    50.616, 50.616, 50.617, 50.617, 50.617, 50.617, 50.618, 50.618, 50.618, 
    50.618, 50.619, 50.619, 50.619, 50.619, 50.62, 50.62, 50.62, 50.62, 
    50.621, 50.621, 50.621, 50.621, 50.622, 50.622, 50.622, 50.622, 50.622, 
    50.623, 50.623, 50.623, 50.623, 50.623, 50.624, 50.624, 50.624, 50.624, 
    50.625, 50.625, 50.625, 50.625, 50.626, 50.626, 50.626, 50.626, 50.626, 
    50.627, 50.627, 50.627, 50.627, 50.628, 50.628, 50.628, 50.629, 50.629, 
    50.629, 50.629, 50.63, 50.63, 50.63, 50.631, 50.631, 50.631, 50.632, 
    50.632, 50.632, 50.632, 50.633, 50.633, 50.633, 50.633, 50.634, 50.634, 
    50.634, 50.635, 50.635, 50.635, 50.635, 50.635, 50.636, 50.636, 50.636, 
    50.636, 50.636, 50.637, 50.637, 50.637, 50.637, 50.638, 50.638, 50.638, 
    50.638, 50.638, 50.639, 50.639, 50.639, 50.639, 50.639, 50.64, 50.64, 
    50.64, 50.64, 50.641, 50.641, 50.641, 50.641, 50.642, 50.642, 50.642, 
    50.642, 50.643, 50.643, 50.643, 50.643, 50.643, 50.644, 50.644, 50.644, 
    50.644, 50.644, 50.645, 50.645, 50.645, 50.645, 50.645, 50.646, 50.646, 
    50.646, 50.646, 50.646, 50.647, 50.647, 50.647, 50.647, 50.648, 50.648, 
    50.648, 50.648, 50.649, 50.649, 50.649, 50.649, 50.65, 50.65, 50.65, 
    50.65, 50.651, 50.651, 50.651, 50.651, 50.651, 50.652, 50.652, 50.652, 
    50.652, 50.653, 50.653, 50.653, 50.653, 50.653, 50.654, 50.654, 50.654, 
    50.654, 50.654, 50.655, 50.655, 50.655, 50.655, 50.655, 50.656, 50.656, 
    50.656, 50.656, 50.657, 50.657, 50.657, 50.657, 50.657, 50.658, 50.658, 
    50.658, 50.658, 50.659, 50.659, 50.659, 50.659, 50.66, 50.66, 50.66, 
    50.66, 50.661, 50.661, 50.661, 50.661, 50.661, 50.662, 50.662, 50.662, 
    50.662, 50.663, 50.663, 50.663, 50.663, 50.663, 50.663, 50.664, 50.664, 
    50.664, 50.664, 50.664, 50.664, 50.665, 50.665, 50.665, 50.665, 50.665, 
    50.665, 50.666, 50.666, 50.666, 50.666, 50.666, 50.666, 50.667, 50.667, 
    50.667, 50.667, 50.667, 50.668, 50.668, 50.668, 50.668, 50.669, 50.669, 
    50.669, 50.669, 50.669, 50.67, 50.67, 50.67, 50.67, 50.671, 50.671, 
    50.671, 50.672, 50.672, 50.672, 50.672, 50.673, 50.673, 50.673, 50.673, 
    50.673, 50.674, 50.674, 50.674, 50.674, 50.675, 50.675, 50.675, 50.675, 
    50.675, 50.676, 50.676, 50.676, 50.676, 50.676, 50.677, 50.677, 50.677, 
    50.677, 50.678, 50.678, 50.678, 50.678, 50.678, 50.679, 50.679, 50.679, 
    50.679, 50.679, 50.68, 50.68, 50.68, 50.68, 50.68, 50.681, 50.681, 
    50.681, 50.681, 50.681, 50.682, 50.682, 50.682, 50.682, 50.682, 50.682, 
    50.683, 50.683, 50.683, 50.683, 50.683, 50.683, 50.684, 50.684, 50.684, 
    50.684, 50.684, 50.685, 50.685, 50.685, 50.685, 50.685, 50.686, 50.686, 
    50.686, 50.686, 50.686, 50.687, 50.687, 50.687, 50.687, 50.687, 50.688, 
    50.688, 50.688, 50.688, 50.688, 50.689, 50.689, 50.689, 50.689, 50.689, 
    50.689, 50.689, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 
    50.691, 50.691, 50.691, 50.691, 50.691, 50.691, 50.691, 50.692, 50.692, 
    50.692, 50.692, 50.692, 50.693, 50.693, 50.693, 50.694, 50.694, 50.694, 
    50.694, 50.695, 50.695, 50.695, 50.696, 50.696, 50.696, 50.697, 50.697, 
    50.697, 50.698, 50.698, 50.698, 50.698, 50.699, 50.699, 50.699, 50.699, 
    50.699, 50.7, 50.7, 50.7, 50.7, 50.7, 50.7, 50.701, 50.701, 50.701, 
    50.701, 50.701, 50.701, 50.701, 50.702, 50.702, 50.702, 50.702, 50.702, 
    50.702, 50.702, 50.703, 50.703, 50.703, 50.703, 50.703, 50.704, 50.704, 
    50.704, 50.704, 50.705, 50.705, 50.705, 50.705, 50.705, 50.706, 50.706, 
    50.706, 50.706, 50.707, 50.707, 50.707, 50.707, 50.707, 50.708, 50.708, 
    50.708, 50.708, 50.709, 50.709, 50.709, 50.709, 50.709, 50.709, 50.71, 
    50.71, 50.71, 50.71, 50.71, 50.71, 50.711, 50.711, 50.711, 50.711, 
    50.711, 50.711, 50.711, 50.711, 50.712, 50.712, 50.712, 50.712, 50.712, 
    50.712, 50.713, 50.713, 50.713, 50.713, 50.714, 50.714, 50.714, 50.714, 
    50.714, 50.715, 50.715, 50.715, 50.715, 50.716, 50.716, 50.716, 50.716, 
    50.716, 50.717, 50.717, 50.717, 50.717, 50.717, 50.717, 50.718, 50.718, 
    50.718, 50.718, 50.718, 50.718, 50.719, 50.719, 50.719, 50.719, 50.719, 
    50.719, 50.72, 50.72, 50.72, 50.72, 50.72, 50.721, 50.721, 50.721, 
    50.721, 50.722, 50.722, 50.722, 50.722, 50.723, 50.723, 50.723, 50.724, 
    50.724, 50.724, 50.724, 50.725, 50.725, 50.725, 50.725, 50.725, 50.726, 
    50.726, 50.726, 50.726, 50.726, 50.726, 50.727, 50.727, 50.727, 50.727, 
    50.727, 50.727, 50.728, 50.728, 50.728, 50.728, 50.728, 50.728, 50.729, 
    50.729, 50.729, 50.729, 50.729, 50.73, 50.73, 50.73, 50.73, 50.73, 
    50.731, 50.731, 50.731, 50.731, 50.731, 50.732, 50.732, 50.732, 50.732, 
    50.732, 50.733, 50.733, 50.733, 50.733, 50.733, 50.734, 50.734, 50.734, 
    50.734, 50.734, 50.734, 50.734, 50.735, 50.735, 50.735, 50.735, 50.735, 
    50.735, 50.735, 50.735, 50.735, 50.736, 50.736, 50.736, 50.736, 50.736, 
    50.736, 50.736, 50.736, 50.737, 50.737, 50.737, 50.737, 50.737, 50.738, 
    50.738, 50.738, 50.738, 50.738, 50.739, 50.739, 50.739, 50.74, 50.74, 
    50.74, 50.74, 50.741, 50.741, 50.741, 50.741, 50.742, 50.742, 50.742, 
    50.742, 50.743, 50.743, 50.743, 50.743, 50.744, 50.744, 50.744, 50.744, 
    50.744, 50.745, 50.745, 50.745, 50.745, 50.745, 50.745, 50.746, 50.746, 
    50.746, 50.746, 50.746, 50.746, 50.746, 50.747, 50.747, 50.747, 50.747, 
    50.747, 50.747, 50.748, 50.748, 50.748, 50.748, 50.748, 50.749, 50.749, 
    50.749, 50.749, 50.75, 50.75, 50.75, 50.751, 50.751, 50.751, 50.751, 
    50.752, 50.752, 50.752, 50.752, 50.752, 50.753, 50.753, 50.753, 50.753, 
    50.754, 50.754, 50.754, 50.754, 50.754, 50.754, 50.755, 50.755, 50.755, 
    50.755, 50.755, 50.755, 50.755, 50.755, 50.756, 50.756, 50.756, 50.756, 
    50.756, 50.756, 50.757, 50.757, 50.757, 50.757, 50.757, 50.757, 50.757, 
    50.758, 50.758, 50.758, 50.758, 50.758, 50.758, 50.758, 50.759, 50.759, 
    50.759, 50.759, 50.759, 50.76, 50.76, 50.76, 50.76, 50.76, 50.76, 50.761, 
    50.761, 50.761, 50.761, 50.762, 50.762, 50.762, 50.762, 50.763, 50.763, 
    50.763, 50.764, 50.764, 50.764, 50.764, 50.765, 50.765, 50.765, 50.765, 
    50.766, 50.766, 50.766, 50.766, 50.766, 50.766, 50.766, 50.767, 50.767, 
    50.767, 50.767, 50.767, 50.767, 50.767, 50.767, 50.768, 50.768, 50.768, 
    50.768, 50.768, 50.768, 50.769, 50.769, 50.769, 50.769, 50.77, 50.77, 
    50.77, 50.77, 50.771, 50.771, 50.771, 50.771, 50.771, 50.772, 50.772, 
    50.772, 50.772, 50.773, 50.773, 50.773, 50.773, 50.773, 50.774, 50.774, 
    50.774, 50.774, 50.774, 50.774, 50.774, 50.775, 50.775, 50.775, 50.775, 
    50.775, 50.775, 50.776, 50.776, 50.776, 50.776, 50.776, 50.777, 50.777, 
    50.777, 50.777, 50.777, 50.778, 50.778, 50.778, 50.778, 50.779, 50.779, 
    50.779, 50.779, 50.779, 50.78, 50.78, 50.78, 50.78, 50.78, 50.78, 50.781, 
    50.781, 50.781, 50.781, 50.781, 50.781, 50.782, 50.782, 50.782, 50.782, 
    50.782, 50.782, 50.783, 50.783, 50.783, 50.783, 50.783, 50.784, 50.784, 
    50.784, 50.784, 50.784, 50.785, 50.785, 50.785, 50.785, 50.785, 50.785, 
    50.786, 50.786, 50.786, 50.786, 50.786, 50.786, 50.787, 50.787, 50.787, 
    50.787, 50.787, 50.787, 50.787, 50.788, 50.788, 50.788, 50.788, 50.788, 
    50.789, 50.789, 50.789, 50.789, 50.79, 50.79, 50.79, 50.79, 50.79, 
    50.791, 50.791, 50.791, 50.791, 50.791, 50.792, 50.792, 50.792, 50.792, 
    50.792, 50.792, 50.793, 50.793, 50.793, 50.793, 50.793, 50.793, 50.793, 
    50.794, 50.794, 50.794, 50.794, 50.794, 50.795, 50.795, 50.795, 50.795, 
    50.796, 50.796, 50.796, 50.796, 50.797, 50.797, 50.797, 50.798, 50.798, 
    50.798, 50.798, 50.799, 50.799, 50.799, 50.799, 50.8, 50.8, 50.8, 50.8, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 50.524, 50.524, 50.525, 50.525, 
    50.525, 50.526, 50.526, 50.527, 50.527, 50.527, 50.528, 50.528, 50.529, 
    50.529, 50.529, 50.53, 50.53, 50.531, 50.531, 50.531, 50.532, 50.532, 
    50.533, 50.533, 50.534, 50.534, 50.535, 50.535, 50.536, 50.536, 50.537, 
    50.537, 50.538, 50.538, 50.539, 50.54, 50.54, 50.541, 50.541, 50.542, 
    50.542, 50.543, 50.543, 50.544, 50.544, 50.544, 50.545, 50.545, 50.546, 
    50.546, 50.546, 50.547, 50.547, 50.547, 50.548, 50.548, 50.548, 50.549, 
    50.549, 50.549, 50.55, 50.55, 50.55, 50.551, 50.551, 50.551, 50.552, 
    50.552, 50.552, 50.553, 50.553, 50.553, 50.554, 50.554, 50.554, 50.555, 
    50.555, 50.555, 50.556, 50.556, 50.556, 50.557, 50.557, 50.557, 50.558, 
    50.558, 50.558, 50.559, 50.559, 50.56, 50.56, 50.56, 50.561, 50.561, 
    50.561, 50.562, 50.562, 50.563, 50.563, 50.563, 50.564, 50.564, 50.565, 
    50.565, 50.565, 50.566, 50.566, 50.567, 50.567, 50.567, 50.568, 50.568, 
    50.568, 50.569, 50.569, 50.57, 50.57, 50.57, 50.571, 50.571, 50.572, 
    50.572, 50.572, 50.573, 50.573, 50.573, 50.574, 50.574, 50.574, 50.575, 
    50.575, 50.575, 50.576, 50.576, 50.576, 50.577, 50.577, 50.577, 50.578, 
    50.578, 50.578, 50.579, 50.579, 50.579, 50.58, 50.58, 50.58, 50.58, 
    50.581, 50.581, 50.581, 50.581, 50.582, 50.582, 50.582, 50.583, 50.583, 
    50.583, 50.584, 50.584, 50.584, 50.584, 50.585, 50.585, 50.585, 50.586, 
    50.586, 50.586, 50.587, 50.587, 50.587, 50.588, 50.588, 50.588, 50.589, 
    50.589, 50.59, 50.59, 50.59, 50.591, 50.591, 50.591, 50.592, 50.592, 
    50.592, 50.593, 50.593, 50.593, 50.594, 50.594, 50.594, 50.595, 50.595, 
    50.595, 50.596, 50.596, 50.596, 50.597, 50.597, 50.597, 50.597, 50.598, 
    50.598, 50.598, 50.598, 50.599, 50.599, 50.599, 50.6, 50.6, 50.6, 50.6, 
    50.601, 50.601, 50.601, 50.602, 50.602, 50.602, 50.603, 50.603, 50.603, 
    50.604, 50.604, 50.604, 50.605, 50.605, 50.605, 50.606, 50.606, 50.606, 
    50.607, 50.607, 50.607, 50.607, 50.608, 50.608, 50.608, 50.608, 50.609, 
    50.609, 50.609, 50.61, 50.61, 50.61, 50.61, 50.61, 50.611, 50.611, 
    50.611, 50.612, 50.612, 50.612, 50.612, 50.613, 50.613, 50.613, 50.613, 
    50.614, 50.614, 50.614, 50.615, 50.615, 50.615, 50.615, 50.616, 50.616, 
    50.616, 50.616, 50.617, 50.617, 50.617, 50.617, 50.618, 50.618, 50.618, 
    50.618, 50.619, 50.619, 50.619, 50.619, 50.62, 50.62, 50.62, 50.62, 
    50.621, 50.621, 50.621, 50.621, 50.622, 50.622, 50.622, 50.622, 50.622, 
    50.623, 50.623, 50.623, 50.623, 50.623, 50.624, 50.624, 50.624, 50.624, 
    50.625, 50.625, 50.625, 50.625, 50.626, 50.626, 50.626, 50.626, 50.626, 
    50.627, 50.627, 50.627, 50.627, 50.628, 50.628, 50.628, 50.629, 50.629, 
    50.629, 50.629, 50.63, 50.63, 50.63, 50.631, 50.631, 50.631, 50.632, 
    50.632, 50.632, 50.632, 50.633, 50.633, 50.633, 50.633, 50.634, 50.634, 
    50.634, 50.635, 50.635, 50.635, 50.635, 50.635, 50.636, 50.636, 50.636, 
    50.636, 50.636, 50.637, 50.637, 50.637, 50.637, 50.638, 50.638, 50.638, 
    50.638, 50.638, 50.639, 50.639, 50.639, 50.639, 50.639, 50.64, 50.64, 
    50.64, 50.64, 50.641, 50.641, 50.641, 50.641, 50.642, 50.642, 50.642, 
    50.642, 50.643, 50.643, 50.643, 50.643, 50.643, 50.644, 50.644, 50.644, 
    50.644, 50.644, 50.645, 50.645, 50.645, 50.645, 50.645, 50.646, 50.646, 
    50.646, 50.646, 50.646, 50.647, 50.647, 50.647, 50.647, 50.648, 50.648, 
    50.648, 50.648, 50.649, 50.649, 50.649, 50.649, 50.65, 50.65, 50.65, 
    50.65, 50.651, 50.651, 50.651, 50.651, 50.651, 50.652, 50.652, 50.652, 
    50.652, 50.653, 50.653, 50.653, 50.653, 50.653, 50.654, 50.654, 50.654, 
    50.654, 50.654, 50.655, 50.655, 50.655, 50.655, 50.655, 50.656, 50.656, 
    50.656, 50.656, 50.657, 50.657, 50.657, 50.657, 50.657, 50.658, 50.658, 
    50.658, 50.658, 50.659, 50.659, 50.659, 50.659, 50.66, 50.66, 50.66, 
    50.66, 50.661, 50.661, 50.661, 50.661, 50.661, 50.662, 50.662, 50.662, 
    50.662, 50.663, 50.663, 50.663, 50.663, 50.663, 50.663, 50.664, 50.664, 
    50.664, 50.664, 50.664, 50.664, 50.665, 50.665, 50.665, 50.665, 50.665, 
    50.665, 50.666, 50.666, 50.666, 50.666, 50.666, 50.666, 50.667, 50.667, 
    50.667, 50.667, 50.667, 50.668, 50.668, 50.668, 50.668, 50.669, 50.669, 
    50.669, 50.669, 50.669, 50.67, 50.67, 50.67, 50.67, 50.671, 50.671, 
    50.671, 50.672, 50.672, 50.672, 50.672, 50.673, 50.673, 50.673, 50.673, 
    50.673, 50.674, 50.674, 50.674, 50.674, 50.675, 50.675, 50.675, 50.675, 
    50.675, 50.676, 50.676, 50.676, 50.676, 50.676, 50.677, 50.677, 50.677, 
    50.677, 50.678, 50.678, 50.678, 50.678, 50.678, 50.679, 50.679, 50.679, 
    50.679, 50.679, 50.68, 50.68, 50.68, 50.68, 50.68, 50.681, 50.681, 
    50.681, 50.681, 50.681, 50.682, 50.682, 50.682, 50.682, 50.682, 50.682, 
    50.683, 50.683, 50.683, 50.683, 50.683, 50.683, 50.684, 50.684, 50.684, 
    50.684, 50.684, 50.685, 50.685, 50.685, 50.685, 50.685, 50.686, 50.686, 
    50.686, 50.686, 50.686, 50.687, 50.687, 50.687, 50.687, 50.687, 50.688, 
    50.688, 50.688, 50.688, 50.688, 50.689, 50.689, 50.689, 50.689, 50.689, 
    50.689, 50.689, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 50.69, 
    50.691, 50.691, 50.691, 50.691, 50.691, 50.691, 50.691, 50.692, 50.692, 
    50.692, 50.692, 50.692, 50.693, 50.693, 50.693, 50.694, 50.694, 50.694, 
    50.694, 50.695, 50.695, 50.695, 50.696, 50.696, 50.696, 50.697, 50.697, 
    50.697, 50.698, 50.698, 50.698, 50.698, 50.699, 50.699, 50.699, 50.699, 
    50.699, 50.7, 50.7, 50.7, 50.7, 50.7, 50.7, 50.701, 50.701, 50.701, 
    50.701, 50.701, 50.701, 50.701, 50.702, 50.702, 50.702, 50.702, 50.702, 
    50.702, 50.702, 50.703, 50.703, 50.703, 50.703, 50.703, 50.704, 50.704, 
    50.704, 50.704, 50.705, 50.705, 50.705, 50.705, 50.705, 50.706, 50.706, 
    50.706, 50.706, 50.707, 50.707, 50.707, 50.707, 50.707, 50.708, 50.708, 
    50.708, 50.708, 50.709, 50.709, 50.709, 50.709, 50.709, 50.709, 50.71, 
    50.71, 50.71, 50.71, 50.71, 50.71, 50.711, 50.711, 50.711, 50.711, 
    50.711, 50.711, 50.711, 50.711, 50.712, 50.712, 50.712, 50.712, 50.712, 
    50.712, 50.713, 50.713, 50.713, 50.713, 50.714, 50.714, 50.714, 50.714, 
    50.714, 50.715, 50.715, 50.715, 50.715, 50.716, 50.716, 50.716, 50.716, 
    50.716, 50.717, 50.717, 50.717, 50.717, 50.717, 50.717, 50.718, 50.718, 
    50.718, 50.718, 50.718, 50.718, 50.719, 50.719, 50.719, 50.719, 50.719, 
    50.719, 50.72, 50.72, 50.72, 50.72, 50.72, 50.721, 50.721, 50.721, 
    50.721, 50.722, 50.722, 50.722, 50.722, 50.723, 50.723, 50.723, 50.724, 
    50.724, 50.724, 50.724, 50.725, 50.725, 50.725, 50.725, 50.725, 50.726, 
    50.726, 50.726, 50.726, 50.726, 50.726, 50.727, 50.727, 50.727, 50.727, 
    50.727, 50.727, 50.728, 50.728, 50.728, 50.728, 50.728, 50.728, 50.729, 
    50.729, 50.729, 50.729, 50.729, 50.73, 50.73, 50.73, 50.73, 50.73, 
    50.731, 50.731, 50.731, 50.731, 50.731, 50.732, 50.732, 50.732, 50.732, 
    50.732, 50.733, 50.733, 50.733, 50.733, 50.733, 50.734, 50.734, 50.734, 
    50.734, 50.734, 50.734, 50.734, 50.735, 50.735, 50.735, 50.735, 50.735, 
    50.735, 50.735, 50.735, 50.735, 50.736, 50.736, 50.736, 50.736, 50.736, 
    50.736, 50.736, 50.736, 50.737, 50.737, 50.737, 50.737, 50.737, 50.738, 
    50.738, 50.738, 50.738, 50.738, 50.739, 50.739, 50.739, 50.74, 50.74, 
    50.74, 50.74, 50.741, 50.741, 50.741, 50.741, 50.742, 50.742, 50.742, 
    50.742, 50.743, 50.743, 50.743, 50.743, 50.744, 50.744, 50.744, 50.744, 
    50.744, 50.745, 50.745, 50.745, 50.745, 50.745, 50.745, 50.746, 50.746, 
    50.746, 50.746, 50.746, 50.746, 50.746, 50.747, 50.747, 50.747, 50.747, 
    50.747, 50.747, 50.748, 50.748, 50.748, 50.748, 50.748, 50.749, 50.749, 
    50.749, 50.749, 50.75, 50.75, 50.75, 50.751, 50.751, 50.751, 50.751, 
    50.752, 50.752, 50.752, 50.752, 50.752, 50.753, 50.753, 50.753, 50.753, 
    50.754, 50.754, 50.754, 50.754, 50.754, 50.754, 50.755, 50.755, 50.755, 
    50.755, 50.755, 50.755, 50.755, 50.755, 50.756, 50.756, 50.756, 50.756, 
    50.756, 50.756, 50.757, 50.757, 50.757, 50.757, 50.757, 50.757, 50.757, 
    50.758, 50.758, 50.758, 50.758, 50.758, 50.758, 50.758, 50.759, 50.759, 
    50.759, 50.759, 50.759, 50.76, 50.76, 50.76, 50.76, 50.76, 50.76, 50.761, 
    50.761, 50.761, 50.761, 50.762, 50.762, 50.762, 50.762, 50.763, 50.763, 
    50.763, 50.764, 50.764, 50.764, 50.764, 50.765, 50.765, 50.765, 50.765, 
    50.766, 50.766, 50.766, 50.766, 50.766, 50.766, 50.766, 50.767, 50.767, 
    50.767, 50.767, 50.767, 50.767, 50.767, 50.767, 50.768, 50.768, 50.768, 
    50.768, 50.768, 50.768, 50.769, 50.769, 50.769, 50.769, 50.77, 50.77, 
    50.77, 50.77, 50.771, 50.771, 50.771, 50.771, 50.771, 50.772, 50.772, 
    50.772, 50.772, 50.773, 50.773, 50.773, 50.773, 50.773, 50.774, 50.774, 
    50.774, 50.774, 50.774, 50.774, 50.774, 50.775, 50.775, 50.775, 50.775, 
    50.775, 50.775, 50.776, 50.776, 50.776, 50.776, 50.776, 50.777, 50.777, 
    50.777, 50.777, 50.777, 50.778, 50.778, 50.778, 50.778, 50.779, 50.779, 
    50.779, 50.779, 50.779, 50.78, 50.78, 50.78, 50.78, 50.78, 50.78, 50.781, 
    50.781, 50.781, 50.781, 50.781, 50.781, 50.782, 50.782, 50.782, 50.782, 
    50.782, 50.782, 50.783, 50.783, 50.783, 50.783, 50.783, 50.784, 50.784, 
    50.784, 50.784, 50.784, 50.785, 50.785, 50.785, 50.785, 50.785, 50.785, 
    50.786, 50.786, 50.786, 50.786, 50.786, 50.786, 50.787, 50.787, 50.787, 
    50.787, 50.787, 50.787, 50.787, 50.788, 50.788, 50.788, 50.788, 50.788, 
    50.789, 50.789, 50.789, 50.789, 50.79, 50.79, 50.79, 50.79, 50.79, 
    50.791, 50.791, 50.791, 50.791, 50.791, 50.792, 50.792, 50.792, 50.792, 
    50.792, 50.792, 50.793, 50.793, 50.793, 50.793, 50.793, 50.793, 50.793, 
    50.794, 50.794, 50.794, 50.794, 50.794, 50.795, 50.795, 50.795, 50.795, 
    50.796, 50.796, 50.796, 50.796, 50.797, 50.797, 50.797, 50.798, 50.798, 
    50.798, 50.798, 50.799, 50.799, 50.799, 50.799, 50.8, 50.8, 50.8, 50.8, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 lon_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -4.015, -4.016, -4.017, -4.017, 
    -4.018, -4.019, -4.019, -4.02, -4.021, -4.021, -4.022, -4.023, -4.023, 
    -4.024, -4.025, -4.025, -4.026, -4.027, -4.027, -4.028, -4.029, -4.029, 
    -4.03, -4.031, -4.031, -4.032, -4.033, -4.033, -4.034, -4.035, -4.035, 
    -4.036, -4.037, -4.037, -4.038, -4.039, -4.039, -4.04, -4.041, -4.041, 
    -4.042, -4.043, -4.043, -4.044, -4.045, -4.045, -4.046, -4.047, -4.047, 
    -4.048, -4.049, -4.049, -4.05, -4.051, -4.051, -4.052, -4.053, -4.053, 
    -4.054, -4.055, -4.055, -4.056, -4.057, -4.057, -4.058, -4.059, -4.06, 
    -4.06, -4.061, -4.062, -4.062, -4.063, -4.064, -4.064, -4.065, -4.066, 
    -4.066, -4.067, -4.068, -4.068, -4.069, -4.07, -4.07, -4.071, -4.072, 
    -4.072, -4.073, -4.074, -4.075, -4.075, -4.076, -4.077, -4.077, -4.078, 
    -4.079, -4.079, -4.08, -4.081, -4.081, -4.082, -4.083, -4.083, -4.084, 
    -4.085, -4.086, -4.086, -4.087, -4.088, -4.088, -4.089, -4.09, -4.09, 
    -4.091, -4.092, -4.092, -4.093, -4.094, -4.094, -4.095, -4.096, -4.096, 
    -4.097, -4.098, -4.098, -4.099, -4.1, -4.101, -4.101, -4.102, -4.103, 
    -4.103, -4.104, -4.105, -4.105, -4.106, -4.107, -4.107, -4.108, -4.109, 
    -4.11, -4.11, -4.111, -4.112, -4.112, -4.113, -4.114, -4.114, -4.115, 
    -4.116, -4.117, -4.117, -4.118, -4.119, -4.119, -4.12, -4.121, -4.122, 
    -4.122, -4.123, -4.124, -4.124, -4.125, -4.126, -4.126, -4.127, -4.128, 
    -4.129, -4.129, -4.13, -4.131, -4.131, -4.132, -4.133, -4.133, -4.134, 
    -4.135, -4.135, -4.136, -4.137, -4.138, -4.138, -4.139, -4.14, -4.14, 
    -4.141, -4.142, -4.142, -4.143, -4.144, -4.144, -4.145, -4.146, -4.147, 
    -4.147, -4.148, -4.149, -4.149, -4.15, -4.151, -4.152, -4.152, -4.153, 
    -4.154, -4.154, -4.155, -4.156, -4.157, -4.157, -4.158, -4.159, -4.159, 
    -4.16, -4.161, -4.162, -4.162, -4.163, -4.164, -4.164, -4.165, -4.166, 
    -4.166, -4.167, -4.168, -4.169, -4.169, -4.17, -4.171, -4.171, -4.172, 
    -4.173, -4.174, -4.174, -4.175, -4.176, -4.176, -4.177, -4.178, -4.179, 
    -4.179, -4.18, -4.181, -4.181, -4.182, -4.183, -4.184, -4.184, -4.185, 
    -4.186, -4.186, -4.187, -4.188, -4.189, -4.189, -4.19, -4.191, -4.192, 
    -4.192, -4.193, -4.194, -4.194, -4.195, -4.196, -4.197, -4.197, -4.198, 
    -4.199, -4.199, -4.2, -4.201, -4.202, -4.202, -4.203, -4.204, -4.204, 
    -4.205, -4.206, -4.207, -4.207, -4.208, -4.209, -4.21, -4.21, -4.211, 
    -4.212, -4.212, -4.213, -4.214, -4.215, -4.215, -4.216, -4.217, -4.218, 
    -4.218, -4.219, -4.22, -4.22, -4.221, -4.222, -4.223, -4.223, -4.224, 
    -4.225, -4.226, -4.226, -4.227, -4.228, -4.229, -4.229, -4.23, -4.231, 
    -4.231, -4.232, -4.233, -4.234, -4.234, -4.235, -4.236, -4.237, -4.237, 
    -4.238, -4.239, -4.239, -4.24, -4.241, -4.242, -4.242, -4.243, -4.244, 
    -4.244, -4.245, -4.246, -4.247, -4.247, -4.248, -4.249, -4.249, -4.25, 
    -4.251, -4.252, -4.252, -4.253, -4.254, -4.255, -4.255, -4.256, -4.257, 
    -4.258, -4.258, -4.259, -4.26, -4.26, -4.261, -4.262, -4.263, -4.263, 
    -4.264, -4.265, -4.266, -4.266, -4.267, -4.268, -4.269, -4.269, -4.27, 
    -4.271, -4.271, -4.272, -4.273, -4.274, -4.274, -4.275, -4.276, -4.277, 
    -4.277, -4.278, -4.279, -4.28, -4.28, -4.281, -4.282, -4.282, -4.283, 
    -4.284, -4.285, -4.285, -4.286, -4.287, -4.288, -4.288, -4.289, -4.29, 
    -4.291, -4.291, -4.292, -4.293, -4.294, -4.294, -4.295, -4.296, -4.297, 
    -4.297, -4.298, -4.299, -4.299, -4.3, -4.301, -4.302, -4.302, -4.303, 
    -4.304, -4.305, -4.305, -4.306, -4.307, -4.307, -4.308, -4.309, -4.31, 
    -4.31, -4.311, -4.312, -4.313, -4.313, -4.314, -4.315, -4.316, -4.316, 
    -4.317, -4.318, -4.319, -4.319, -4.32, -4.321, -4.322, -4.322, -4.323, 
    -4.324, -4.324, -4.325, -4.326, -4.327, -4.327, -4.328, -4.329, -4.33, 
    -4.33, -4.331, -4.332, -4.333, -4.333, -4.334, -4.335, -4.335, -4.336, 
    -4.337, -4.338, -4.338, -4.339, -4.34, -4.341, -4.341, -4.342, -4.343, 
    -4.344, -4.344, -4.345, -4.346, -4.347, -4.347, -4.348, -4.349, -4.35, 
    -4.35, -4.351, -4.352, -4.352, -4.353, -4.354, -4.355, -4.355, -4.356, 
    -4.357, -4.358, -4.358, -4.359, -4.36, -4.361, -4.361, -4.362, -4.363, 
    -4.364, -4.364, -4.365, -4.366, -4.367, -4.367, -4.368, -4.369, -4.37, 
    -4.37, -4.371, -4.372, -4.373, -4.373, -4.374, -4.375, -4.375, -4.376, 
    -4.377, -4.378, -4.378, -4.379, -4.38, -4.381, -4.381, -4.382, -4.383, 
    -4.384, -4.384, -4.385, -4.386, -4.387, -4.387, -4.388, -4.389, -4.389, 
    -4.39, -4.391, -4.392, -4.392, -4.393, -4.394, -4.395, -4.395, -4.396, 
    -4.397, -4.398, -4.398, -4.399, -4.4, -4.401, -4.401, -4.402, -4.403, 
    -4.404, -4.404, -4.405, -4.406, -4.406, -4.407, -4.408, -4.409, -4.409, 
    -4.41, -4.411, -4.412, -4.412, -4.413, -4.414, -4.415, -4.415, -4.416, 
    -4.417, -4.418, -4.418, -4.419, -4.42, -4.421, -4.421, -4.422, -4.423, 
    -4.424, -4.424, -4.425, -4.426, -4.427, -4.427, -4.428, -4.429, -4.43, 
    -4.43, -4.431, -4.432, -4.433, -4.433, -4.434, -4.435, -4.435, -4.436, 
    -4.437, -4.438, -4.438, -4.439, -4.44, -4.441, -4.441, -4.442, -4.443, 
    -4.444, -4.444, -4.445, -4.446, -4.447, -4.447, -4.448, -4.449, -4.45, 
    -4.45, -4.451, -4.452, -4.453, -4.453, -4.454, -4.455, -4.456, -4.456, 
    -4.457, -4.458, -4.459, -4.459, -4.46, -4.461, -4.462, -4.462, -4.463, 
    -4.464, -4.465, -4.465, -4.466, -4.467, -4.467, -4.468, -4.469, -4.47, 
    -4.47, -4.471, -4.472, -4.473, -4.473, -4.474, -4.475, -4.475, -4.476, 
    -4.477, -4.478, -4.478, -4.479, -4.48, -4.481, -4.481, -4.482, -4.483, 
    -4.484, -4.484, -4.485, -4.486, -4.487, -4.487, -4.488, -4.489, -4.49, 
    -4.49, -4.491, -4.492, -4.493, -4.493, -4.494, -4.495, -4.496, -4.496, 
    -4.497, -4.498, -4.499, -4.499, -4.5, -4.501, -4.502, -4.502, -4.503, 
    -4.504, -4.504, -4.505, -4.506, -4.507, -4.507, -4.508, -4.509, -4.51, 
    -4.51, -4.511, -4.512, -4.513, -4.513, -4.514, -4.515, -4.516, -4.516, 
    -4.517, -4.518, -4.519, -4.519, -4.52, -4.521, -4.522, -4.522, -4.523, 
    -4.524, -4.525, -4.525, -4.526, -4.527, -4.528, -4.528, -4.529, -4.53, 
    -4.531, -4.531, -4.532, -4.533, -4.534, -4.534, -4.535, -4.536, -4.536, 
    -4.537, -4.538, -4.539, -4.539, -4.54, -4.541, -4.542, -4.542, -4.543, 
    -4.544, -4.545, -4.545, -4.546, -4.547, -4.548, -4.548, -4.549, -4.55, 
    -4.551, -4.551, -4.552, -4.553, -4.554, -4.554, -4.555, -4.556, -4.557, 
    -4.557, -4.558, -4.559, -4.559, -4.56, -4.561, -4.562, -4.562, -4.563, 
    -4.564, -4.565, -4.565, -4.566, -4.567, -4.568, -4.568, -4.569, -4.57, 
    -4.571, -4.571, -4.572, -4.573, -4.573, -4.574, -4.575, -4.576, -4.576, 
    -4.577, -4.578, -4.579, -4.579, -4.58, -4.581, -4.582, -4.582, -4.583, 
    -4.584, -4.585, -4.585, -4.586, -4.587, -4.588, -4.588, -4.589, -4.59, 
    -4.591, -4.591, -4.592, -4.593, -4.594, -4.594, -4.595, -4.596, -4.596, 
    -4.597, -4.598, -4.599, -4.599, -4.6, -4.601, -4.602, -4.602, -4.603, 
    -4.604, -4.605, -4.605, -4.606, -4.607, -4.608, -4.608, -4.609, -4.61, 
    -4.611, -4.611, -4.612, -4.613, -4.614, -4.614, -4.615, -4.616, -4.617, 
    -4.617, -4.618, -4.619, -4.62, -4.62, -4.621, -4.622, -4.623, -4.623, 
    -4.624, -4.625, -4.626, -4.626, -4.627, -4.628, -4.629, -4.629, -4.63, 
    -4.631, -4.632, -4.632, -4.633, -4.634, -4.635, -4.635, -4.636, -4.637, 
    -4.637, -4.638, -4.639, -4.64, -4.64, -4.641, -4.642, -4.643, -4.643, 
    -4.644, -4.645, -4.645, -4.646, -4.647, -4.648, -4.648, -4.649, -4.65, 
    -4.651, -4.651, -4.652, -4.653, -4.654, -4.654, -4.655, -4.656, -4.657, 
    -4.657, -4.658, -4.659, -4.66, -4.66, -4.661, -4.662, -4.663, -4.663, 
    -4.664, -4.665, -4.666, -4.666, -4.667, -4.668, -4.669, -4.669, -4.67, 
    -4.671, -4.671, -4.672, -4.673, -4.674, -4.674, -4.675, -4.676, -4.677, 
    -4.677, -4.678, -4.679, -4.679, -4.68, -4.681, -4.682, -4.682, -4.683, 
    -4.684, -4.685, -4.685, -4.686, -4.687, -4.688, -4.688, -4.689, -4.69, 
    -4.691, -4.691, -4.692, -4.693, -4.694, -4.694, -4.695, -4.696, -4.697, 
    -4.697, -4.698, -4.699, -4.7, -4.7, -4.701, -4.702, -4.703, -4.703, 
    -4.704, -4.705, -4.706, -4.706, -4.707, -4.708, -4.709, -4.709, -4.71, 
    -4.711, -4.711, -4.712, -4.713, -4.714, -4.714, -4.715, -4.716, -4.717, 
    -4.717, -4.718, -4.719, -4.72, -4.72, -4.721, -4.722, -4.723, -4.723, 
    -4.724, -4.725, -4.726, -4.726, -4.727, -4.728, -4.728, -4.729, -4.73, 
    -4.731, -4.731, -4.732, -4.733, -4.734, -4.734, -4.735, -4.736, -4.737, 
    -4.737, -4.738, -4.739, -4.74, -4.74, -4.741, -4.742, -4.743, -4.743, 
    -4.744, -4.745, -4.746, -4.746, -4.747, -4.748, -4.748, -4.749, -4.75, 
    -4.751, -4.751, -4.752, -4.753, -4.754, -4.754, -4.755, -4.756, -4.757, 
    -4.757, -4.758, -4.759, -4.76, -4.76, -4.761, -4.762, -4.762, -4.763, 
    -4.764, -4.765, -4.765, -4.766, -4.767, -4.768, -4.768, -4.769, -4.77, 
    -4.771, -4.771, -4.772, -4.773, -4.774, -4.774, -4.775, -4.776, -4.777, 
    -4.777, -4.778, -4.779, -4.78, -4.78, -4.781, -4.782, -4.782, -4.783, 
    -4.784, -4.785, -4.785, -4.786, -4.787, -4.788, -4.788, -4.789, -4.79, 
    -4.791, -4.791, -4.792, -4.793, -4.794, -4.794, -4.795, -4.796, -4.797, 
    -4.797, -4.798, -4.799, -4.8, -4.8, -4.801, -4.802, -4.802, -4.803, 
    -4.804, -4.805, -4.805, -4.806, -4.807, -4.808, -4.808, -4.809, -4.81, 
    -4.811, -4.811, -4.812, -4.813, -4.814, -4.814, -4.815, -4.816, -4.817, 
    -4.817, -4.818, -4.819, -4.82, -4.82, -4.821, -4.822, -4.822, -4.823, 
    -4.824, -4.825, -4.825, -4.826, -4.827, -4.828, -4.828, -4.829, -4.83, 
    -4.831, -4.831, -4.832, -4.833, -4.834, -4.834, -4.835, -4.836, -4.836, 
    -4.837, -4.838, -4.839, -4.839, -4.84, -4.841, -4.842, -4.842, -4.843, 
    -4.844, -4.845, -4.845, -4.846, -4.847, -4.848, -4.848, -4.849, -4.85, 
    -4.851, -4.851, -4.852, -4.853, -4.854, -4.854, -4.855, -4.856, -4.856, 
    -4.857, -4.858, -4.859, -4.859, -4.86, -4.861, -4.862, -4.862, -4.863, 
    -4.864, -4.864, -4.865, -4.866, -4.867, -4.867, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -4.015, -4.016, -4.017, -4.017, 
    -4.018, -4.019, -4.019, -4.02, -4.021, -4.021, -4.022, -4.023, -4.023, 
    -4.024, -4.025, -4.025, -4.026, -4.027, -4.027, -4.028, -4.029, -4.029, 
    -4.03, -4.031, -4.031, -4.032, -4.033, -4.033, -4.034, -4.035, -4.035, 
    -4.036, -4.037, -4.037, -4.038, -4.039, -4.039, -4.04, -4.041, -4.041, 
    -4.042, -4.043, -4.043, -4.044, -4.045, -4.045, -4.046, -4.047, -4.047, 
    -4.048, -4.049, -4.049, -4.05, -4.051, -4.051, -4.052, -4.053, -4.053, 
    -4.054, -4.055, -4.055, -4.056, -4.057, -4.057, -4.058, -4.059, -4.06, 
    -4.06, -4.061, -4.062, -4.062, -4.063, -4.064, -4.064, -4.065, -4.066, 
    -4.066, -4.067, -4.068, -4.068, -4.069, -4.07, -4.07, -4.071, -4.072, 
    -4.072, -4.073, -4.074, -4.075, -4.075, -4.076, -4.077, -4.077, -4.078, 
    -4.079, -4.079, -4.08, -4.081, -4.081, -4.082, -4.083, -4.083, -4.084, 
    -4.085, -4.086, -4.086, -4.087, -4.088, -4.088, -4.089, -4.09, -4.09, 
    -4.091, -4.092, -4.092, -4.093, -4.094, -4.094, -4.095, -4.096, -4.096, 
    -4.097, -4.098, -4.098, -4.099, -4.1, -4.101, -4.101, -4.102, -4.103, 
    -4.103, -4.104, -4.105, -4.105, -4.106, -4.107, -4.107, -4.108, -4.109, 
    -4.11, -4.11, -4.111, -4.112, -4.112, -4.113, -4.114, -4.114, -4.115, 
    -4.116, -4.117, -4.117, -4.118, -4.119, -4.119, -4.12, -4.121, -4.122, 
    -4.122, -4.123, -4.124, -4.124, -4.125, -4.126, -4.126, -4.127, -4.128, 
    -4.129, -4.129, -4.13, -4.131, -4.131, -4.132, -4.133, -4.133, -4.134, 
    -4.135, -4.135, -4.136, -4.137, -4.138, -4.138, -4.139, -4.14, -4.14, 
    -4.141, -4.142, -4.142, -4.143, -4.144, -4.144, -4.145, -4.146, -4.147, 
    -4.147, -4.148, -4.149, -4.149, -4.15, -4.151, -4.152, -4.152, -4.153, 
    -4.154, -4.154, -4.155, -4.156, -4.157, -4.157, -4.158, -4.159, -4.159, 
    -4.16, -4.161, -4.162, -4.162, -4.163, -4.164, -4.164, -4.165, -4.166, 
    -4.166, -4.167, -4.168, -4.169, -4.169, -4.17, -4.171, -4.171, -4.172, 
    -4.173, -4.174, -4.174, -4.175, -4.176, -4.176, -4.177, -4.178, -4.179, 
    -4.179, -4.18, -4.181, -4.181, -4.182, -4.183, -4.184, -4.184, -4.185, 
    -4.186, -4.186, -4.187, -4.188, -4.189, -4.189, -4.19, -4.191, -4.192, 
    -4.192, -4.193, -4.194, -4.194, -4.195, -4.196, -4.197, -4.197, -4.198, 
    -4.199, -4.199, -4.2, -4.201, -4.202, -4.202, -4.203, -4.204, -4.204, 
    -4.205, -4.206, -4.207, -4.207, -4.208, -4.209, -4.21, -4.21, -4.211, 
    -4.212, -4.212, -4.213, -4.214, -4.215, -4.215, -4.216, -4.217, -4.218, 
    -4.218, -4.219, -4.22, -4.22, -4.221, -4.222, -4.223, -4.223, -4.224, 
    -4.225, -4.226, -4.226, -4.227, -4.228, -4.229, -4.229, -4.23, -4.231, 
    -4.231, -4.232, -4.233, -4.234, -4.234, -4.235, -4.236, -4.237, -4.237, 
    -4.238, -4.239, -4.239, -4.24, -4.241, -4.242, -4.242, -4.243, -4.244, 
    -4.244, -4.245, -4.246, -4.247, -4.247, -4.248, -4.249, -4.249, -4.25, 
    -4.251, -4.252, -4.252, -4.253, -4.254, -4.255, -4.255, -4.256, -4.257, 
    -4.258, -4.258, -4.259, -4.26, -4.26, -4.261, -4.262, -4.263, -4.263, 
    -4.264, -4.265, -4.266, -4.266, -4.267, -4.268, -4.269, -4.269, -4.27, 
    -4.271, -4.271, -4.272, -4.273, -4.274, -4.274, -4.275, -4.276, -4.277, 
    -4.277, -4.278, -4.279, -4.28, -4.28, -4.281, -4.282, -4.282, -4.283, 
    -4.284, -4.285, -4.285, -4.286, -4.287, -4.288, -4.288, -4.289, -4.29, 
    -4.291, -4.291, -4.292, -4.293, -4.294, -4.294, -4.295, -4.296, -4.297, 
    -4.297, -4.298, -4.299, -4.299, -4.3, -4.301, -4.302, -4.302, -4.303, 
    -4.304, -4.305, -4.305, -4.306, -4.307, -4.307, -4.308, -4.309, -4.31, 
    -4.31, -4.311, -4.312, -4.313, -4.313, -4.314, -4.315, -4.316, -4.316, 
    -4.317, -4.318, -4.319, -4.319, -4.32, -4.321, -4.322, -4.322, -4.323, 
    -4.324, -4.324, -4.325, -4.326, -4.327, -4.327, -4.328, -4.329, -4.33, 
    -4.33, -4.331, -4.332, -4.333, -4.333, -4.334, -4.335, -4.335, -4.336, 
    -4.337, -4.338, -4.338, -4.339, -4.34, -4.341, -4.341, -4.342, -4.343, 
    -4.344, -4.344, -4.345, -4.346, -4.347, -4.347, -4.348, -4.349, -4.35, 
    -4.35, -4.351, -4.352, -4.352, -4.353, -4.354, -4.355, -4.355, -4.356, 
    -4.357, -4.358, -4.358, -4.359, -4.36, -4.361, -4.361, -4.362, -4.363, 
    -4.364, -4.364, -4.365, -4.366, -4.367, -4.367, -4.368, -4.369, -4.37, 
    -4.37, -4.371, -4.372, -4.373, -4.373, -4.374, -4.375, -4.375, -4.376, 
    -4.377, -4.378, -4.378, -4.379, -4.38, -4.381, -4.381, -4.382, -4.383, 
    -4.384, -4.384, -4.385, -4.386, -4.387, -4.387, -4.388, -4.389, -4.389, 
    -4.39, -4.391, -4.392, -4.392, -4.393, -4.394, -4.395, -4.395, -4.396, 
    -4.397, -4.398, -4.398, -4.399, -4.4, -4.401, -4.401, -4.402, -4.403, 
    -4.404, -4.404, -4.405, -4.406, -4.406, -4.407, -4.408, -4.409, -4.409, 
    -4.41, -4.411, -4.412, -4.412, -4.413, -4.414, -4.415, -4.415, -4.416, 
    -4.417, -4.418, -4.418, -4.419, -4.42, -4.421, -4.421, -4.422, -4.423, 
    -4.424, -4.424, -4.425, -4.426, -4.427, -4.427, -4.428, -4.429, -4.43, 
    -4.43, -4.431, -4.432, -4.433, -4.433, -4.434, -4.435, -4.435, -4.436, 
    -4.437, -4.438, -4.438, -4.439, -4.44, -4.441, -4.441, -4.442, -4.443, 
    -4.444, -4.444, -4.445, -4.446, -4.447, -4.447, -4.448, -4.449, -4.45, 
    -4.45, -4.451, -4.452, -4.453, -4.453, -4.454, -4.455, -4.456, -4.456, 
    -4.457, -4.458, -4.459, -4.459, -4.46, -4.461, -4.462, -4.462, -4.463, 
    -4.464, -4.465, -4.465, -4.466, -4.467, -4.467, -4.468, -4.469, -4.47, 
    -4.47, -4.471, -4.472, -4.473, -4.473, -4.474, -4.475, -4.475, -4.476, 
    -4.477, -4.478, -4.478, -4.479, -4.48, -4.481, -4.481, -4.482, -4.483, 
    -4.484, -4.484, -4.485, -4.486, -4.487, -4.487, -4.488, -4.489, -4.49, 
    -4.49, -4.491, -4.492, -4.493, -4.493, -4.494, -4.495, -4.496, -4.496, 
    -4.497, -4.498, -4.499, -4.499, -4.5, -4.501, -4.502, -4.502, -4.503, 
    -4.504, -4.504, -4.505, -4.506, -4.507, -4.507, -4.508, -4.509, -4.51, 
    -4.51, -4.511, -4.512, -4.513, -4.513, -4.514, -4.515, -4.516, -4.516, 
    -4.517, -4.518, -4.519, -4.519, -4.52, -4.521, -4.522, -4.522, -4.523, 
    -4.524, -4.525, -4.525, -4.526, -4.527, -4.528, -4.528, -4.529, -4.53, 
    -4.531, -4.531, -4.532, -4.533, -4.534, -4.534, -4.535, -4.536, -4.536, 
    -4.537, -4.538, -4.539, -4.539, -4.54, -4.541, -4.542, -4.542, -4.543, 
    -4.544, -4.545, -4.545, -4.546, -4.547, -4.548, -4.548, -4.549, -4.55, 
    -4.551, -4.551, -4.552, -4.553, -4.554, -4.554, -4.555, -4.556, -4.557, 
    -4.557, -4.558, -4.559, -4.559, -4.56, -4.561, -4.562, -4.562, -4.563, 
    -4.564, -4.565, -4.565, -4.566, -4.567, -4.568, -4.568, -4.569, -4.57, 
    -4.571, -4.571, -4.572, -4.573, -4.573, -4.574, -4.575, -4.576, -4.576, 
    -4.577, -4.578, -4.579, -4.579, -4.58, -4.581, -4.582, -4.582, -4.583, 
    -4.584, -4.585, -4.585, -4.586, -4.587, -4.588, -4.588, -4.589, -4.59, 
    -4.591, -4.591, -4.592, -4.593, -4.594, -4.594, -4.595, -4.596, -4.596, 
    -4.597, -4.598, -4.599, -4.599, -4.6, -4.601, -4.602, -4.602, -4.603, 
    -4.604, -4.605, -4.605, -4.606, -4.607, -4.608, -4.608, -4.609, -4.61, 
    -4.611, -4.611, -4.612, -4.613, -4.614, -4.614, -4.615, -4.616, -4.617, 
    -4.617, -4.618, -4.619, -4.62, -4.62, -4.621, -4.622, -4.623, -4.623, 
    -4.624, -4.625, -4.626, -4.626, -4.627, -4.628, -4.629, -4.629, -4.63, 
    -4.631, -4.632, -4.632, -4.633, -4.634, -4.635, -4.635, -4.636, -4.637, 
    -4.637, -4.638, -4.639, -4.64, -4.64, -4.641, -4.642, -4.643, -4.643, 
    -4.644, -4.645, -4.645, -4.646, -4.647, -4.648, -4.648, -4.649, -4.65, 
    -4.651, -4.651, -4.652, -4.653, -4.654, -4.654, -4.655, -4.656, -4.657, 
    -4.657, -4.658, -4.659, -4.66, -4.66, -4.661, -4.662, -4.663, -4.663, 
    -4.664, -4.665, -4.666, -4.666, -4.667, -4.668, -4.669, -4.669, -4.67, 
    -4.671, -4.671, -4.672, -4.673, -4.674, -4.674, -4.675, -4.676, -4.677, 
    -4.677, -4.678, -4.679, -4.679, -4.68, -4.681, -4.682, -4.682, -4.683, 
    -4.684, -4.685, -4.685, -4.686, -4.687, -4.688, -4.688, -4.689, -4.69, 
    -4.691, -4.691, -4.692, -4.693, -4.694, -4.694, -4.695, -4.696, -4.697, 
    -4.697, -4.698, -4.699, -4.7, -4.7, -4.701, -4.702, -4.703, -4.703, 
    -4.704, -4.705, -4.706, -4.706, -4.707, -4.708, -4.709, -4.709, -4.71, 
    -4.711, -4.711, -4.712, -4.713, -4.714, -4.714, -4.715, -4.716, -4.717, 
    -4.717, -4.718, -4.719, -4.72, -4.72, -4.721, -4.722, -4.723, -4.723, 
    -4.724, -4.725, -4.726, -4.726, -4.727, -4.728, -4.728, -4.729, -4.73, 
    -4.731, -4.731, -4.732, -4.733, -4.734, -4.734, -4.735, -4.736, -4.737, 
    -4.737, -4.738, -4.739, -4.74, -4.74, -4.741, -4.742, -4.743, -4.743, 
    -4.744, -4.745, -4.746, -4.746, -4.747, -4.748, -4.748, -4.749, -4.75, 
    -4.751, -4.751, -4.752, -4.753, -4.754, -4.754, -4.755, -4.756, -4.757, 
    -4.757, -4.758, -4.759, -4.76, -4.76, -4.761, -4.762, -4.762, -4.763, 
    -4.764, -4.765, -4.765, -4.766, -4.767, -4.768, -4.768, -4.769, -4.77, 
    -4.771, -4.771, -4.772, -4.773, -4.774, -4.774, -4.775, -4.776, -4.777, 
    -4.777, -4.778, -4.779, -4.78, -4.78, -4.781, -4.782, -4.782, -4.783, 
    -4.784, -4.785, -4.785, -4.786, -4.787, -4.788, -4.788, -4.789, -4.79, 
    -4.791, -4.791, -4.792, -4.793, -4.794, -4.794, -4.795, -4.796, -4.797, 
    -4.797, -4.798, -4.799, -4.8, -4.8, -4.801, -4.802, -4.802, -4.803, 
    -4.804, -4.805, -4.805, -4.806, -4.807, -4.808, -4.808, -4.809, -4.81, 
    -4.811, -4.811, -4.812, -4.813, -4.814, -4.814, -4.815, -4.816, -4.817, 
    -4.817, -4.818, -4.819, -4.82, -4.82, -4.821, -4.822, -4.822, -4.823, 
    -4.824, -4.825, -4.825, -4.826, -4.827, -4.828, -4.828, -4.829, -4.83, 
    -4.831, -4.831, -4.832, -4.833, -4.834, -4.834, -4.835, -4.836, -4.836, 
    -4.837, -4.838, -4.839, -4.839, -4.84, -4.841, -4.842, -4.842, -4.843, 
    -4.844, -4.845, -4.845, -4.846, -4.847, -4.848, -4.848, -4.849, -4.85, 
    -4.851, -4.851, -4.852, -4.853, -4.854, -4.854, -4.855, -4.856, -4.856, 
    -4.857, -4.858, -4.859, -4.859, -4.86, -4.861, -4.862, -4.862, -4.863, 
    -4.864, -4.864, -4.865, -4.866, -4.867, -4.867, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 azimuth_tp =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 193.13, 193.13, 193.13, 193.13, 
    193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 
    193.13, 193.13, 193.13, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 
    193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 
    193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.11, 193.11, 193.11, 
    193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 
    193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.1, 193.1, 
    193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 
    193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.09, 193.09, 193.09, 
    193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 
    193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.08, 193.08, 
    193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 
    193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 
    193.08, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 
    193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 
    193.07, 193.07, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 
    193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 
    193.06, 193.06, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 
    193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 
    193.05, 193.05, 193.05, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 
    193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 
    193.04, 193.04, 193.04, 193.04, 193.04, 193.03, 193.03, 193.03, 193.03, 
    193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 
    193.03, 193.03, 193.03, 193.03, 193.03, 193.02, 193.02, 193.02, 193.02, 
    193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 
    193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.01, 193.01, 193.01, 
    193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 
    193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193, 193, 193, 193, 193, 
    193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 
    192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 
    192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 
    192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 
    192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 
    192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 
    192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 
    192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 
    192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 
    192.96, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 
    192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 
    192.95, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 
    192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 
    192.94, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 
    192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 
    192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 
    192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 
    192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 
    192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 
    192.91, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 
    192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.89, 
    192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 
    192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.88, 192.88, 
    192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 
    192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.87, 192.87, 
    192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 
    192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.86, 192.86, 192.86, 
    192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 
    192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.85, 192.85, 
    192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 
    192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.84, 192.84, 
    192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 
    192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.83, 192.83, 
    192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 
    192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.82, 192.82, 192.82, 
    192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 
    192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.81, 192.81, 192.81, 
    192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 
    192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.8, 192.8, 192.8, 
    192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 
    192.8, 192.8, 192.8, 192.8, 192.8, 192.79, 192.79, 192.79, 192.79, 
    192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 
    192.79, 192.79, 192.79, 192.79, 192.79, 192.78, 192.78, 192.78, 192.78, 
    192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 
    192.78, 192.78, 192.78, 192.78, 192.77, 192.77, 192.77, 192.77, 192.77, 
    192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 
    192.77, 192.77, 192.77, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 
    192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 
    192.76, 192.76, 192.76, 192.76, 192.75, 192.75, 192.75, 192.75, 192.75, 
    192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 
    192.75, 192.75, 192.75, 192.75, 192.74, 192.74, 192.74, 192.74, 192.74, 
    192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 
    192.74, 192.74, 192.74, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 
    192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 
    192.73, 192.73, 192.73, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 
    192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 
    192.72, 192.72, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 
    192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 
    192.71, 192.71, 192.71, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 
    192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 
    192.7, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 
    192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 
    192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 
    192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 
    192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 
    192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.66, 
    192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 
    192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.65, 
    192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 
    192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 
    192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 
    192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.63, 
    192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 
    192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.62, 
    192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 
    192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.61, 192.61, 
    192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 
    192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.6, 192.6, 
    192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 
    192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.59, 192.59, 192.59, 
    192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 
    192.59, 192.59, 192.59, 192.59, 192.59, 192.58, 192.58, 192.58, 192.58, 
    192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 
    192.58, 192.58, 192.58, 192.58, 192.58, 192.57, 192.57, 192.57, 192.57, 
    192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 
    192.57, 192.57, 192.57, 192.57, 192.57, 192.56, 192.56, 192.56, 192.56, 
    192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 
    192.56, 192.56, 192.56, 192.56, 192.55, 192.55, 192.55, 192.55, 192.55, 
    192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 
    192.55, 192.55, 192.55, 192.55, 192.54, 192.54, 192.54, 192.54, 192.54, 
    192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 
    192.54, 192.54, 192.54, 192.54, 192.54, 192.53, 192.53, 192.53, 192.53, 
    192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 
    192.53, 192.53, 192.53, 192.53, 192.52, 192.52, 192.52, 192.52, 192.52, 
    192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 
    192.52, 192.52, 192.52, 192.52, 192.51, 192.51, 192.51, 192.51, 192.51, 
    192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 
    192.51, 192.51, 192.51, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 
    192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 
    192.5, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 
    192.49, 192.49, 192.49, 192.49, 192.49, 192.49, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 193.13, 193.13, 193.13, 193.13, 
    193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 193.13, 
    193.13, 193.13, 193.13, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 
    193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 
    193.12, 193.12, 193.12, 193.12, 193.12, 193.12, 193.11, 193.11, 193.11, 
    193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 
    193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.11, 193.1, 193.1, 
    193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 
    193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.1, 193.09, 193.09, 193.09, 
    193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 
    193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.09, 193.08, 193.08, 
    193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 
    193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 193.08, 
    193.08, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 
    193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 193.07, 
    193.07, 193.07, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 
    193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 193.06, 
    193.06, 193.06, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 
    193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 193.05, 
    193.05, 193.05, 193.05, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 
    193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 193.04, 
    193.04, 193.04, 193.04, 193.04, 193.04, 193.03, 193.03, 193.03, 193.03, 
    193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 193.03, 
    193.03, 193.03, 193.03, 193.03, 193.03, 193.02, 193.02, 193.02, 193.02, 
    193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 
    193.02, 193.02, 193.02, 193.02, 193.02, 193.02, 193.01, 193.01, 193.01, 
    193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 
    193.01, 193.01, 193.01, 193.01, 193.01, 193.01, 193, 193, 193, 193, 193, 
    193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 
    192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 
    192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 192.99, 
    192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 
    192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 192.98, 
    192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 
    192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 192.97, 
    192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 
    192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 192.96, 
    192.96, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 
    192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 192.95, 
    192.95, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 
    192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 192.94, 
    192.94, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 
    192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 192.93, 
    192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 
    192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 192.92, 
    192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 
    192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 192.91, 
    192.91, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 
    192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.9, 192.89, 
    192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 
    192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.89, 192.88, 192.88, 
    192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 
    192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.88, 192.87, 192.87, 
    192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 
    192.87, 192.87, 192.87, 192.87, 192.87, 192.87, 192.86, 192.86, 192.86, 
    192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 
    192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.86, 192.85, 192.85, 
    192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 
    192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.85, 192.84, 192.84, 
    192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 
    192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.84, 192.83, 192.83, 
    192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 
    192.83, 192.83, 192.83, 192.83, 192.83, 192.83, 192.82, 192.82, 192.82, 
    192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 
    192.82, 192.82, 192.82, 192.82, 192.82, 192.82, 192.81, 192.81, 192.81, 
    192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 
    192.81, 192.81, 192.81, 192.81, 192.81, 192.81, 192.8, 192.8, 192.8, 
    192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 192.8, 
    192.8, 192.8, 192.8, 192.8, 192.8, 192.79, 192.79, 192.79, 192.79, 
    192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 192.79, 
    192.79, 192.79, 192.79, 192.79, 192.79, 192.78, 192.78, 192.78, 192.78, 
    192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 192.78, 
    192.78, 192.78, 192.78, 192.78, 192.77, 192.77, 192.77, 192.77, 192.77, 
    192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 192.77, 
    192.77, 192.77, 192.77, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 
    192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 192.76, 
    192.76, 192.76, 192.76, 192.76, 192.75, 192.75, 192.75, 192.75, 192.75, 
    192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 192.75, 
    192.75, 192.75, 192.75, 192.75, 192.74, 192.74, 192.74, 192.74, 192.74, 
    192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 192.74, 
    192.74, 192.74, 192.74, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 
    192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 192.73, 
    192.73, 192.73, 192.73, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 
    192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 192.72, 
    192.72, 192.72, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 
    192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 192.71, 
    192.71, 192.71, 192.71, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 
    192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 192.7, 
    192.7, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 
    192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 192.69, 
    192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 
    192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 192.68, 
    192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 
    192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.67, 192.66, 
    192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 
    192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.66, 192.65, 
    192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 
    192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 192.65, 
    192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 
    192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.64, 192.63, 
    192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 
    192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.63, 192.62, 
    192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 
    192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.62, 192.61, 192.61, 
    192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 
    192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.61, 192.6, 192.6, 
    192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 
    192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.6, 192.59, 192.59, 192.59, 
    192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 192.59, 
    192.59, 192.59, 192.59, 192.59, 192.59, 192.58, 192.58, 192.58, 192.58, 
    192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 192.58, 
    192.58, 192.58, 192.58, 192.58, 192.58, 192.57, 192.57, 192.57, 192.57, 
    192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 192.57, 
    192.57, 192.57, 192.57, 192.57, 192.57, 192.56, 192.56, 192.56, 192.56, 
    192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 192.56, 
    192.56, 192.56, 192.56, 192.56, 192.55, 192.55, 192.55, 192.55, 192.55, 
    192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 192.55, 
    192.55, 192.55, 192.55, 192.55, 192.54, 192.54, 192.54, 192.54, 192.54, 
    192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 192.54, 
    192.54, 192.54, 192.54, 192.54, 192.54, 192.53, 192.53, 192.53, 192.53, 
    192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 192.53, 
    192.53, 192.53, 192.53, 192.53, 192.52, 192.52, 192.52, 192.52, 192.52, 
    192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 192.52, 
    192.52, 192.52, 192.52, 192.52, 192.51, 192.51, 192.51, 192.51, 192.51, 
    192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 192.51, 
    192.51, 192.51, 192.51, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 
    192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 192.5, 
    192.5, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 192.49, 
    192.49, 192.49, 192.49, 192.49, 192.49, 192.49, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 impact_L1 =
  6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.377e+06, 6.377e+06, 
    6.377e+06, 6.377e+06, 6.3771e+06, 6.3771e+06, 6.3772e+06, 6.3772e+06, 
    6.3772e+06, 6.3773e+06, 6.3773e+06, 6.3774e+06, 6.3774e+06, 6.3775e+06, 
    6.3775e+06, 6.3775e+06, 6.3776e+06, 6.3776e+06, 6.3777e+06, 6.3777e+06, 
    6.3777e+06, 6.3777e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3782e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 
    6.3784e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3786e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.3789e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3786e+06, 6.3786e+06, 6.3786e+06, 
    6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3784e+06, 
    6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 
    6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3782e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3781e+06, 6.3781e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 6.3784e+06, 
    6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3796e+06, 
    6.3796e+06, 6.3796e+06, 6.3797e+06, 6.3797e+06, 6.3798e+06, 6.3798e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.38e+06, 
    6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3798e+06, 6.3798e+06, 
    6.3798e+06, 6.3798e+06, 6.3797e+06, 6.3797e+06, 6.3796e+06, 6.3796e+06, 
    6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3794e+06, 6.3794e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3805e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3805e+06, 6.3805e+06, 
    6.3805e+06, 6.3805e+06, 6.3805e+06, 6.3806e+06, 6.3806e+06, 6.3806e+06, 
    6.3807e+06, 6.3807e+06, 6.3807e+06, 6.3808e+06, 6.3808e+06, 6.3808e+06, 
    6.3809e+06, 6.3809e+06, 6.3809e+06, 6.381e+06, 6.381e+06, 6.381e+06, 
    6.381e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 
    6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 
    6.3815e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 
    6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 
    6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 
    6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 
    6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 
    6.382e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 
    6.3821e+06, 6.3821e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 
    6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3823e+06, 6.3823e+06, 
    6.3823e+06, 6.3823e+06, 6.3823e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 
    6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3825e+06, 6.3825e+06, 
    6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 
    6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3827e+06, 
    6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3828e+06, 6.3828e+06, 
    6.3828e+06, 6.3828e+06, 6.3828e+06, 6.3829e+06, 6.3829e+06, 6.3829e+06, 
    6.3829e+06, 6.3829e+06, 6.383e+06, 6.383e+06, 6.383e+06, 6.383e+06, 
    6.383e+06, 6.383e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 
    6.3831e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 
    6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 
    6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3837e+06, 
    6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3838e+06, 
    6.3838e+06, 6.3838e+06, 6.3838e+06, 6.3839e+06, 6.3839e+06, 6.3839e+06, 
    6.3839e+06, 6.3839e+06, 6.3839e+06, 6.384e+06, 6.384e+06, 6.384e+06, 
    6.384e+06, 6.384e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 
    6.3841e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3843e+06, 
    6.3843e+06, 6.3843e+06, 6.3843e+06, 6.3844e+06, 6.3844e+06, 6.3844e+06, 
    6.3844e+06, 6.3845e+06, 6.3845e+06, 6.3845e+06, 6.3846e+06, 6.3846e+06, 
    6.3846e+06, 6.3846e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 
    6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3849e+06, 
    6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.385e+06, 
    6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 
    6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 
    6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3853e+06, 
    6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3854e+06, 
    6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3855e+06, 6.3855e+06, 
    6.3855e+06, 6.3855e+06, 6.3855e+06, 6.3856e+06, 6.3856e+06, 6.3856e+06, 
    6.3856e+06, 6.3856e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 
    6.3857e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3859e+06, 
    6.3859e+06, 6.3859e+06, 6.3859e+06, 6.3859e+06, 6.386e+06, 6.386e+06, 
    6.386e+06, 6.386e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.3951e+06, 6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3962e+06, 6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 
    6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3975e+06, 6.3975e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 
    6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 
    6.3983e+06, 6.3983e+06, 6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3986e+06, 6.3986e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3993e+06, 6.3993e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3995e+06, 
    6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 
    6.4006e+06, 6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 
    6.4008e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 
    6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 
    6.4017e+06, 6.4017e+06, 6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 
    6.4029e+06, 6.4029e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4037e+06, 
    6.4037e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 
    6.404e+06, 6.4041e+06, 6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 
    6.405e+06, 6.405e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 
    6.406e+06, 6.406e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 
    6.4063e+06, 6.4063e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 6.4065e+06, 
    6.4066e+06, 6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 
    6.4069e+06, 6.4069e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4072e+06, 6.4072e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4079e+06, 6.4079e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4082e+06, 6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 6.4084e+06, 
    6.4085e+06, 6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4088e+06, 
    6.4088e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.4091e+06, 
    6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4095e+06, 6.4095e+06, 6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 
    6.4098e+06, 6.4099e+06, 6.4099e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 
    6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4107e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 6.411e+06, 6.4111e+06, 
    6.4111e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 
    6.4115e+06, 6.4115e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4119e+06, 6.4119e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 
    6.4121e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4124e+06, 
    6.4125e+06, 6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4128e+06, 
    6.4128e+06, 6.4129e+06, 6.4129e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 6.4138e+06, 
    6.4138e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.4141e+06, 
    6.4141e+06, 6.4142e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 
    6.4148e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.4151e+06, 6.4151e+06, 
    6.4152e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4155e+06, 
    6.4156e+06, 6.4156e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4159e+06, 
    6.4159e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 6.4161e+06, 6.4162e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 6.4165e+06, 
    6.4166e+06, 6.4166e+06, 6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 6.4172e+06, 
    6.4172e+06, 6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 
    6.4179e+06, 6.418e+06, 6.418e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 
    6.4183e+06, 6.4183e+06, 6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 6.4189e+06, 
    6.419e+06, 6.419e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 6.42e+06, 
    6.42e+06, 6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 
    6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 6.4206e+06, 6.4207e+06, 
    6.4207e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 
    6.4211e+06, 6.4211e+06, 6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 6.4217e+06, 
    6.4218e+06, 6.4218e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.4221e+06, 
    6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 6.4227e+06, 6.4228e+06, 
    6.4229e+06, 6.4229e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 6.4232e+06, 
    6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 6.4238e+06, 
    6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 6.4241e+06, 6.4241e+06, 
    6.4242e+06, 6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4245e+06, 
    6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 6.4252e+06, 
    6.4252e+06, 6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4258e+06, 6.4258e+06, 6.4259e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 6.4262e+06, 
    6.4263e+06, 6.4264e+06, 6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 
    6.4266e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 
    6.427e+06, 6.427e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 
    6.4277e+06, 6.4277e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 6.4283e+06, 6.4283e+06, 
    6.4284e+06, 6.4284e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4287e+06, 
    6.4288e+06, 6.4288e+06, 6.4289e+06, 6.4289e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 6.4294e+06, 
    6.4295e+06, 6.4295e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.43e+06, 6.43e+06, 6.4301e+06, 
    6.4301e+06, 6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 6.4312e+06, 
    6.4312e+06, 6.4313e+06, 6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4318e+06, 6.4318e+06, 
    6.4319e+06, 6.4319e+06, 6.432e+06, 6.432e+06, 6.4321e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 
    6.4326e+06, 6.4326e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 6.4331e+06, 6.4332e+06, 
    6.4333e+06, 6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4336e+06, 
    6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4343e+06, 
    6.4343e+06, 6.4344e+06, 6.4344e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 6.4349e+06, 
    6.435e+06, 6.4351e+06, 6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 
    6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4356e+06, 6.4357e+06, 
    6.4357e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 6.436e+06, 
    6.4361e+06, 6.4362e+06, 6.4362e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 
    6.4368e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 6.4371e+06, 
    6.4372e+06, 6.4372e+06, 6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 
    6.4375e+06, 6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4378e+06, 
    6.4378e+06, 6.4379e+06, 6.4379e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4384e+06, 
    6.4385e+06, 6.4386e+06, 6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.4391e+06, 6.4392e+06, 
    6.4392e+06, 6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4395e+06, 6.4395e+06, 
    6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 
    6.4399e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4402e+06, 
    6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 
    6.4406e+06, 6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4409e+06, 
    6.4409e+06, 6.441e+06, 6.441e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 6.4416e+06, 
    6.4416e+06, 6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.4421e+06, 6.4421e+06, 6.4422e+06, 6.4422e+06, 6.4423e+06, 
    6.4423e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4427e+06, 6.4428e+06, 6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4433e+06, 6.4434e+06, 
    6.4434e+06, 6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 6.444e+06, 6.444e+06, 
    6.4441e+06, 6.4441e+06, 6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 
    6.4444e+06, 6.4445e+06, 6.4445e+06, 6.4446e+06, 6.4446e+06, 6.4447e+06, 
    6.4447e+06, 6.4448e+06, 6.4449e+06, 6.4449e+06, 6.445e+06, 6.445e+06, 
    6.4451e+06, 6.4452e+06, 6.4452e+06, 6.4453e+06, 6.4453e+06, 6.4454e+06, 
    6.4455e+06, 6.4455e+06, 6.4456e+06, 6.4457e+06, 6.4457e+06, 6.4458e+06, 
    6.4458e+06, 6.4459e+06, 6.4459e+06, 6.446e+06, 6.4461e+06, 6.4461e+06, 
    6.4462e+06, 6.4462e+06, 6.4463e+06, 6.4463e+06, 6.4464e+06, 6.4465e+06, 
    6.4465e+06, 6.4466e+06, 6.4466e+06, 6.4467e+06, 6.4467e+06, 6.4468e+06, 
    6.4468e+06, 6.4469e+06, 6.447e+06, 6.447e+06, 6.4471e+06, 6.4471e+06, 
    6.4472e+06, 6.4472e+06, 6.4473e+06, 6.4474e+06, 6.4474e+06, 6.4475e+06, 
    6.4475e+06, 6.4476e+06, 6.4477e+06, 6.4477e+06, 6.4478e+06, 6.4478e+06, 
    6.4479e+06, 6.448e+06, 6.448e+06, 6.4481e+06, 6.4481e+06, 6.4482e+06, 
    6.4482e+06, 6.4483e+06, 6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4485e+06, 
    6.4486e+06, 6.4486e+06, 6.4487e+06, 6.4487e+06, 6.4488e+06, 6.4489e+06, 
    6.4489e+06, 6.449e+06, 6.449e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 
    6.4493e+06, 6.4493e+06, 6.4494e+06, 6.4494e+06, 6.4495e+06, 6.4496e+06, 
    6.4496e+06, 6.4497e+06, 6.4497e+06, 6.4498e+06, 6.4499e+06, 6.4499e+06, 
    6.45e+06, 6.45e+06, 6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 
    6.4503e+06, 6.4504e+06, 6.4504e+06, 6.4505e+06, 6.4506e+06, 6.4506e+06, 
    6.4507e+06, 6.4507e+06, 6.4508e+06, 6.4508e+06, 6.4509e+06, 6.451e+06, 
    6.451e+06, 6.4511e+06, 6.4511e+06, 6.4512e+06, 6.4513e+06, 6.4513e+06, 
    6.4514e+06, 6.4514e+06, 6.4515e+06, 6.4516e+06, 6.4516e+06, 6.4517e+06, 
    6.4517e+06, 6.4518e+06, 6.4518e+06, 6.4519e+06, 6.452e+06, 6.452e+06, 
    6.4521e+06, 6.4521e+06, 6.4522e+06, 6.4522e+06, 6.4523e+06, 6.4524e+06, 
    6.4524e+06, 6.4525e+06, 6.4525e+06, 6.4526e+06, 6.4526e+06, 6.4527e+06, 
    6.4527e+06, 6.4528e+06, 6.4529e+06, 6.4529e+06, 6.453e+06, 6.453e+06, 
    6.4531e+06, 6.4532e+06, 6.4532e+06, 6.4533e+06, 6.4533e+06, 6.4534e+06, 
    6.4535e+06, 6.4535e+06, 6.4536e+06, 6.4536e+06, 6.4537e+06, 6.4538e+06, 
    6.4538e+06, 6.4539e+06, 6.4539e+06, 6.454e+06, 6.454e+06, 6.4541e+06, 
    6.4541e+06, 6.4542e+06, 6.4543e+06, 6.4543e+06, 6.4544e+06, 6.4544e+06, 
    6.4545e+06, 6.4545e+06, 6.4546e+06, 6.4546e+06, 6.4547e+06, 6.4547e+06, 
    6.4548e+06, 6.4548e+06, 6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 
    6.4551e+06, 6.4552e+06, 6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 
    6.4555e+06, 6.4555e+06, 6.4556e+06, 6.4557e+06, 6.4557e+06, 6.4558e+06, 
    6.4559e+06, 6.4559e+06, 6.456e+06, 6.456e+06, 6.4561e+06, 6.4562e+06, 
    6.4562e+06, 6.4563e+06, 6.4563e+06, 6.4564e+06, 6.4565e+06, 6.4565e+06, 
    6.4566e+06, 6.4566e+06, 6.4567e+06, 6.4567e+06, 6.4568e+06, 6.4568e+06, 
    6.4569e+06,
  6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.377e+06, 6.377e+06, 
    6.377e+06, 6.377e+06, 6.3771e+06, 6.3771e+06, 6.3772e+06, 6.3772e+06, 
    6.3772e+06, 6.3773e+06, 6.3773e+06, 6.3774e+06, 6.3774e+06, 6.3775e+06, 
    6.3775e+06, 6.3775e+06, 6.3776e+06, 6.3776e+06, 6.3777e+06, 6.3777e+06, 
    6.3777e+06, 6.3777e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3782e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 
    6.3784e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3786e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.3789e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3786e+06, 6.3786e+06, 6.3786e+06, 
    6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3784e+06, 
    6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 
    6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3782e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3781e+06, 6.3781e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 6.3784e+06, 
    6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3796e+06, 
    6.3796e+06, 6.3796e+06, 6.3797e+06, 6.3797e+06, 6.3798e+06, 6.3798e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.38e+06, 
    6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3798e+06, 6.3798e+06, 
    6.3798e+06, 6.3798e+06, 6.3797e+06, 6.3797e+06, 6.3796e+06, 6.3796e+06, 
    6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3794e+06, 6.3794e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3805e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3805e+06, 6.3805e+06, 
    6.3805e+06, 6.3805e+06, 6.3805e+06, 6.3806e+06, 6.3806e+06, 6.3806e+06, 
    6.3807e+06, 6.3807e+06, 6.3807e+06, 6.3808e+06, 6.3808e+06, 6.3808e+06, 
    6.3809e+06, 6.3809e+06, 6.3809e+06, 6.381e+06, 6.381e+06, 6.381e+06, 
    6.381e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 
    6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 
    6.3815e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 
    6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 
    6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 
    6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 
    6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 
    6.382e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 
    6.3821e+06, 6.3821e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 
    6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3823e+06, 6.3823e+06, 
    6.3823e+06, 6.3823e+06, 6.3823e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 
    6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3825e+06, 6.3825e+06, 
    6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 
    6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3827e+06, 
    6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3828e+06, 6.3828e+06, 
    6.3828e+06, 6.3828e+06, 6.3828e+06, 6.3829e+06, 6.3829e+06, 6.3829e+06, 
    6.3829e+06, 6.3829e+06, 6.383e+06, 6.383e+06, 6.383e+06, 6.383e+06, 
    6.383e+06, 6.383e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 
    6.3831e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 
    6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 
    6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3837e+06, 
    6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3838e+06, 
    6.3838e+06, 6.3838e+06, 6.3838e+06, 6.3839e+06, 6.3839e+06, 6.3839e+06, 
    6.3839e+06, 6.3839e+06, 6.3839e+06, 6.384e+06, 6.384e+06, 6.384e+06, 
    6.384e+06, 6.384e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 
    6.3841e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3843e+06, 
    6.3843e+06, 6.3843e+06, 6.3843e+06, 6.3844e+06, 6.3844e+06, 6.3844e+06, 
    6.3844e+06, 6.3845e+06, 6.3845e+06, 6.3845e+06, 6.3846e+06, 6.3846e+06, 
    6.3846e+06, 6.3846e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 
    6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3849e+06, 
    6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.385e+06, 
    6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 
    6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 
    6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3853e+06, 
    6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3854e+06, 
    6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3855e+06, 6.3855e+06, 
    6.3855e+06, 6.3855e+06, 6.3855e+06, 6.3856e+06, 6.3856e+06, 6.3856e+06, 
    6.3856e+06, 6.3856e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 
    6.3857e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3859e+06, 
    6.3859e+06, 6.3859e+06, 6.3859e+06, 6.3859e+06, 6.386e+06, 6.386e+06, 
    6.386e+06, 6.386e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.3951e+06, 6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3962e+06, 6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 
    6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3975e+06, 6.3975e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 
    6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 
    6.3983e+06, 6.3983e+06, 6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3986e+06, 6.3986e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3993e+06, 6.3993e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3995e+06, 
    6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 
    6.4006e+06, 6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 
    6.4008e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 
    6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 
    6.4017e+06, 6.4017e+06, 6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 
    6.4029e+06, 6.4029e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4037e+06, 
    6.4037e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 
    6.404e+06, 6.4041e+06, 6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 
    6.405e+06, 6.405e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 
    6.406e+06, 6.406e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 
    6.4063e+06, 6.4063e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 6.4065e+06, 
    6.4066e+06, 6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 
    6.4069e+06, 6.4069e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4072e+06, 6.4072e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4079e+06, 6.4079e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4082e+06, 6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 6.4084e+06, 
    6.4085e+06, 6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4088e+06, 
    6.4088e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.4091e+06, 
    6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4095e+06, 6.4095e+06, 6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 
    6.4098e+06, 6.4099e+06, 6.4099e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 
    6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4107e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 6.411e+06, 6.4111e+06, 
    6.4111e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 
    6.4115e+06, 6.4115e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4119e+06, 6.4119e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 
    6.4121e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4124e+06, 
    6.4125e+06, 6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4128e+06, 
    6.4128e+06, 6.4129e+06, 6.4129e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 6.4138e+06, 
    6.4138e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.4141e+06, 
    6.4141e+06, 6.4142e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 
    6.4148e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.4151e+06, 6.4151e+06, 
    6.4152e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4155e+06, 
    6.4156e+06, 6.4156e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4159e+06, 
    6.4159e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 6.4161e+06, 6.4162e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 6.4165e+06, 
    6.4166e+06, 6.4166e+06, 6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 6.4172e+06, 
    6.4172e+06, 6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 
    6.4179e+06, 6.418e+06, 6.418e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 
    6.4183e+06, 6.4183e+06, 6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 6.4189e+06, 
    6.419e+06, 6.419e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 6.42e+06, 
    6.42e+06, 6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 
    6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 6.4206e+06, 6.4207e+06, 
    6.4207e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 
    6.4211e+06, 6.4211e+06, 6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 6.4217e+06, 
    6.4218e+06, 6.4218e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.4221e+06, 
    6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 6.4227e+06, 6.4228e+06, 
    6.4229e+06, 6.4229e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 6.4232e+06, 
    6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 6.4238e+06, 
    6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 6.4241e+06, 6.4241e+06, 
    6.4242e+06, 6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4245e+06, 
    6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 6.4252e+06, 
    6.4252e+06, 6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4258e+06, 6.4258e+06, 6.4259e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 6.4262e+06, 
    6.4263e+06, 6.4264e+06, 6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 
    6.4266e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 
    6.427e+06, 6.427e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 
    6.4277e+06, 6.4277e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 6.4283e+06, 6.4283e+06, 
    6.4284e+06, 6.4284e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4287e+06, 
    6.4288e+06, 6.4288e+06, 6.4289e+06, 6.4289e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 6.4294e+06, 
    6.4295e+06, 6.4295e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.43e+06, 6.43e+06, 6.4301e+06, 
    6.4301e+06, 6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 6.4312e+06, 
    6.4312e+06, 6.4313e+06, 6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4318e+06, 6.4318e+06, 
    6.4319e+06, 6.4319e+06, 6.432e+06, 6.432e+06, 6.4321e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 
    6.4326e+06, 6.4326e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 6.4331e+06, 6.4332e+06, 
    6.4333e+06, 6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4336e+06, 
    6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4343e+06, 
    6.4343e+06, 6.4344e+06, 6.4344e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 6.4349e+06, 
    6.435e+06, 6.4351e+06, 6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 
    6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4356e+06, 6.4357e+06, 
    6.4357e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 6.436e+06, 
    6.4361e+06, 6.4362e+06, 6.4362e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 
    6.4368e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 6.4371e+06, 
    6.4372e+06, 6.4372e+06, 6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 
    6.4375e+06, 6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4378e+06, 
    6.4378e+06, 6.4379e+06, 6.4379e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4384e+06, 
    6.4385e+06, 6.4386e+06, 6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.4391e+06, 6.4392e+06, 
    6.4392e+06, 6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4395e+06, 6.4395e+06, 
    6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 
    6.4399e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4402e+06, 
    6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 
    6.4406e+06, 6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4409e+06, 
    6.4409e+06, 6.441e+06, 6.441e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 6.4416e+06, 
    6.4416e+06, 6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.4421e+06, 6.4421e+06, 6.4422e+06, 6.4422e+06, 6.4423e+06, 
    6.4423e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4427e+06, 6.4428e+06, 6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4433e+06, 6.4434e+06, 
    6.4434e+06, 6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 6.444e+06, 6.444e+06, 
    6.4441e+06, 6.4441e+06, 6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 
    6.4444e+06, 6.4445e+06, 6.4445e+06, 6.4446e+06, 6.4446e+06, 6.4447e+06, 
    6.4447e+06, 6.4448e+06, 6.4449e+06, 6.4449e+06, 6.445e+06, 6.445e+06, 
    6.4451e+06, 6.4452e+06, 6.4452e+06, 6.4453e+06, 6.4453e+06, 6.4454e+06, 
    6.4455e+06, 6.4455e+06, 6.4456e+06, 6.4457e+06, 6.4457e+06, 6.4458e+06, 
    6.4458e+06, 6.4459e+06, 6.4459e+06, 6.446e+06, 6.4461e+06, 6.4461e+06, 
    6.4462e+06, 6.4462e+06, 6.4463e+06, 6.4463e+06, 6.4464e+06, 6.4465e+06, 
    6.4465e+06, 6.4466e+06, 6.4466e+06, 6.4467e+06, 6.4467e+06, 6.4468e+06, 
    6.4468e+06, 6.4469e+06, 6.447e+06, 6.447e+06, 6.4471e+06, 6.4471e+06, 
    6.4472e+06, 6.4472e+06, 6.4473e+06, 6.4474e+06, 6.4474e+06, 6.4475e+06, 
    6.4475e+06, 6.4476e+06, 6.4477e+06, 6.4477e+06, 6.4478e+06, 6.4478e+06, 
    6.4479e+06, 6.448e+06, 6.448e+06, 6.4481e+06, 6.4481e+06, 6.4482e+06, 
    6.4482e+06, 6.4483e+06, 6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4485e+06, 
    6.4486e+06, 6.4486e+06, 6.4487e+06, 6.4487e+06, 6.4488e+06, 6.4489e+06, 
    6.4489e+06, 6.449e+06, 6.449e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 
    6.4493e+06, 6.4493e+06, 6.4494e+06, 6.4494e+06, 6.4495e+06, 6.4496e+06, 
    6.4496e+06, 6.4497e+06, 6.4497e+06, 6.4498e+06, 6.4499e+06, 6.4499e+06, 
    6.45e+06, 6.45e+06, 6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 
    6.4503e+06, 6.4504e+06, 6.4504e+06, 6.4505e+06, 6.4506e+06, 6.4506e+06, 
    6.4507e+06, 6.4507e+06, 6.4508e+06, 6.4508e+06, 6.4509e+06, 6.451e+06, 
    6.451e+06, 6.4511e+06, 6.4511e+06, 6.4512e+06, 6.4513e+06, 6.4513e+06, 
    6.4514e+06, 6.4514e+06, 6.4515e+06, 6.4516e+06, 6.4516e+06, 6.4517e+06, 
    6.4517e+06, 6.4518e+06, 6.4518e+06, 6.4519e+06, 6.452e+06, 6.452e+06, 
    6.4521e+06, 6.4521e+06, 6.4522e+06, 6.4522e+06, 6.4523e+06, 6.4524e+06, 
    6.4524e+06, 6.4525e+06, 6.4525e+06, 6.4526e+06, 6.4526e+06, 6.4527e+06, 
    6.4527e+06, 6.4528e+06, 6.4529e+06, 6.4529e+06, 6.453e+06, 6.453e+06, 
    6.4531e+06, 6.4532e+06, 6.4532e+06, 6.4533e+06, 6.4533e+06, 6.4534e+06, 
    6.4535e+06, 6.4535e+06, 6.4536e+06, 6.4536e+06, 6.4537e+06, 6.4538e+06, 
    6.4538e+06, 6.4539e+06, 6.4539e+06, 6.454e+06, 6.454e+06, 6.4541e+06, 
    6.4541e+06, 6.4542e+06, 6.4543e+06, 6.4543e+06, 6.4544e+06, 6.4544e+06, 
    6.4545e+06, 6.4545e+06, 6.4546e+06, 6.4546e+06, 6.4547e+06, 6.4547e+06, 
    6.4548e+06, 6.4548e+06, 6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 
    6.4551e+06, 6.4552e+06, 6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 
    6.4555e+06, 6.4555e+06, 6.4556e+06, 6.4557e+06, 6.4557e+06, 6.4558e+06, 
    6.4559e+06, 6.4559e+06, 6.456e+06, 6.456e+06, 6.4561e+06, 6.4562e+06, 
    6.4562e+06, 6.4563e+06, 6.4563e+06, 6.4564e+06, 6.4565e+06, 6.4565e+06, 
    6.4566e+06, 6.4566e+06, 6.4567e+06, 6.4567e+06, 6.4568e+06, 6.4568e+06, 
    6.4569e+06 ;

 impact_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 6.3946e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 6.3955e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3962e+06, 6.3962e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 6.3968e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3976e+06, 6.3976e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3978e+06, 
    6.3978e+06, 6.3979e+06, 6.3979e+06, 6.398e+06, 6.398e+06, 6.3981e+06, 
    6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 6.3983e+06, 6.3983e+06, 
    6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 6.3986e+06, 6.3986e+06, 
    6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 6.3988e+06, 6.3989e+06, 
    6.3989e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.3991e+06, 6.3991e+06, 
    6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3993e+06, 6.3993e+06, 6.3994e+06, 
    6.3994e+06, 6.3994e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3996e+06, 
    6.3996e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3998e+06, 6.3998e+06, 
    6.3999e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 6.4e+06, 6.4001e+06, 
    6.4001e+06, 6.4002e+06, 6.4002e+06, 6.4003e+06, 6.4003e+06, 6.4004e+06, 
    6.4004e+06, 6.4005e+06, 6.4005e+06, 6.4005e+06, 6.4006e+06, 6.4006e+06, 
    6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 6.4009e+06, 6.4009e+06, 
    6.401e+06, 6.401e+06, 6.4011e+06, 6.4011e+06, 6.4011e+06, 6.4012e+06, 
    6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4014e+06, 6.4014e+06, 6.4015e+06, 
    6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 6.4017e+06, 6.4017e+06, 
    6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 6.402e+06, 6.402e+06, 
    6.4021e+06, 6.4021e+06, 6.4022e+06, 6.4022e+06, 6.4023e+06, 6.4023e+06, 
    6.4024e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 6.4026e+06, 6.4026e+06, 
    6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 6.4029e+06, 6.4029e+06, 
    6.403e+06, 6.403e+06, 6.4031e+06, 6.4031e+06, 6.4032e+06, 6.4032e+06, 
    6.4033e+06, 6.4033e+06, 6.4034e+06, 6.4034e+06, 6.4035e+06, 6.4035e+06, 
    6.4036e+06, 6.4036e+06, 6.4037e+06, 6.4037e+06, 6.4038e+06, 6.4038e+06, 
    6.4039e+06, 6.4039e+06, 6.404e+06, 6.404e+06, 6.4041e+06, 6.4041e+06, 
    6.4042e+06, 6.4042e+06, 6.4043e+06, 6.4043e+06, 6.4044e+06, 6.4044e+06, 
    6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 6.4047e+06, 6.4048e+06, 
    6.4048e+06, 6.4049e+06, 6.4049e+06, 6.405e+06, 6.405e+06, 6.4051e+06, 
    6.4051e+06, 6.4052e+06, 6.4052e+06, 6.4053e+06, 6.4054e+06, 6.4054e+06, 
    6.4055e+06, 6.4055e+06, 6.4056e+06, 6.4056e+06, 6.4057e+06, 6.4057e+06, 
    6.4058e+06, 6.4058e+06, 6.4059e+06, 6.406e+06, 6.406e+06, 6.4061e+06, 
    6.4061e+06, 6.4062e+06, 6.4062e+06, 6.4063e+06, 6.4063e+06, 6.4064e+06, 
    6.4064e+06, 6.4065e+06, 6.4065e+06, 6.4065e+06, 6.4066e+06, 6.4066e+06, 
    6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 6.4069e+06, 6.4069e+06, 
    6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 6.4072e+06, 6.4072e+06, 
    6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 6.4075e+06, 6.4076e+06, 
    6.4076e+06, 6.4077e+06, 6.4077e+06, 6.4078e+06, 6.4078e+06, 6.4079e+06, 
    6.408e+06, 6.408e+06, 6.4081e+06, 6.4081e+06, 6.4082e+06, 6.4082e+06, 
    6.4083e+06, 6.4084e+06, 6.4084e+06, 6.4085e+06, 6.4085e+06, 6.4086e+06, 
    6.4086e+06, 6.4087e+06, 6.4087e+06, 6.4088e+06, 6.4088e+06, 6.4089e+06, 
    6.409e+06, 6.409e+06, 6.4091e+06, 6.4091e+06, 6.4092e+06, 6.4092e+06, 
    6.4093e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 6.4095e+06, 6.4096e+06, 
    6.4096e+06, 6.4097e+06, 6.4097e+06, 6.4098e+06, 6.4098e+06, 6.4099e+06, 
    6.41e+06, 6.41e+06, 6.4101e+06, 6.4101e+06, 6.4102e+06, 6.4102e+06, 
    6.4103e+06, 6.4104e+06, 6.4104e+06, 6.4105e+06, 6.4105e+06, 6.4106e+06, 
    6.4106e+06, 6.4107e+06, 6.4107e+06, 6.4108e+06, 6.4108e+06, 6.4109e+06, 
    6.411e+06, 6.411e+06, 6.4111e+06, 6.4111e+06, 6.4112e+06, 6.4112e+06, 
    6.4113e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 6.4115e+06, 6.4115e+06, 
    6.4116e+06, 6.4117e+06, 6.4117e+06, 6.4118e+06, 6.4118e+06, 6.4119e+06, 
    6.4119e+06, 6.412e+06, 6.4121e+06, 6.4121e+06, 6.4122e+06, 6.4122e+06, 
    6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4125e+06, 6.4125e+06, 6.4126e+06, 
    6.4126e+06, 6.4127e+06, 6.4127e+06, 6.4128e+06, 6.4129e+06, 6.4129e+06, 
    6.413e+06, 6.413e+06, 6.4131e+06, 6.4131e+06, 6.4132e+06, 6.4132e+06, 
    6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 6.4135e+06, 6.4136e+06, 
    6.4136e+06, 6.4137e+06, 6.4137e+06, 6.4138e+06, 6.4138e+06, 6.4139e+06, 
    6.4139e+06, 6.414e+06, 6.4141e+06, 6.4141e+06, 6.4142e+06, 6.4142e+06, 
    6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4145e+06, 6.4145e+06, 6.4146e+06, 
    6.4146e+06, 6.4147e+06, 6.4148e+06, 6.4148e+06, 6.4149e+06, 6.4149e+06, 
    6.415e+06, 6.4151e+06, 6.4151e+06, 6.4152e+06, 6.4152e+06, 6.4153e+06, 
    6.4154e+06, 6.4154e+06, 6.4155e+06, 6.4156e+06, 6.4156e+06, 6.4157e+06, 
    6.4157e+06, 6.4158e+06, 6.4158e+06, 6.4159e+06, 6.416e+06, 6.416e+06, 
    6.4161e+06, 6.4161e+06, 6.4162e+06, 6.4162e+06, 6.4163e+06, 6.4164e+06, 
    6.4164e+06, 6.4165e+06, 6.4165e+06, 6.4166e+06, 6.4166e+06, 6.4167e+06, 
    6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 6.4169e+06, 6.417e+06, 
    6.4171e+06, 6.4171e+06, 6.4172e+06, 6.4172e+06, 6.4173e+06, 6.4173e+06, 
    6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 6.4176e+06, 6.4177e+06, 
    6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 6.4179e+06, 6.418e+06, 
    6.4181e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 6.4183e+06, 6.4183e+06, 
    6.4184e+06, 6.4185e+06, 6.4185e+06, 6.4186e+06, 6.4186e+06, 6.4187e+06, 
    6.4187e+06, 6.4188e+06, 6.4189e+06, 6.4189e+06, 6.419e+06, 6.419e+06, 
    6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4193e+06, 6.4193e+06, 6.4194e+06, 
    6.4194e+06, 6.4195e+06, 6.4196e+06, 6.4196e+06, 6.4197e+06, 6.4197e+06, 
    6.4198e+06, 6.4199e+06, 6.4199e+06, 6.42e+06, 6.42e+06, 6.4201e+06, 
    6.4202e+06, 6.4202e+06, 6.4203e+06, 6.4203e+06, 6.4204e+06, 6.4205e+06, 
    6.4205e+06, 6.4206e+06, 6.4206e+06, 6.4207e+06, 6.4207e+06, 6.4208e+06, 
    6.4209e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 6.4211e+06, 6.4212e+06, 
    6.4212e+06, 6.4213e+06, 6.4213e+06, 6.4214e+06, 6.4214e+06, 6.4215e+06, 
    6.4216e+06, 6.4216e+06, 6.4217e+06, 6.4217e+06, 6.4218e+06, 6.4219e+06, 
    6.4219e+06, 6.422e+06, 6.422e+06, 6.4221e+06, 6.4222e+06, 6.4222e+06, 
    6.4223e+06, 6.4224e+06, 6.4224e+06, 6.4225e+06, 6.4226e+06, 6.4226e+06, 
    6.4227e+06, 6.4228e+06, 6.4228e+06, 6.4229e+06, 6.4229e+06, 6.423e+06, 
    6.4231e+06, 6.4231e+06, 6.4232e+06, 6.4232e+06, 6.4233e+06, 6.4234e+06, 
    6.4234e+06, 6.4235e+06, 6.4235e+06, 6.4236e+06, 6.4236e+06, 6.4237e+06, 
    6.4237e+06, 6.4238e+06, 6.4238e+06, 6.4239e+06, 6.4239e+06, 6.424e+06, 
    6.424e+06, 6.4241e+06, 6.4241e+06, 6.4242e+06, 6.4242e+06, 6.4243e+06, 
    6.4243e+06, 6.4244e+06, 6.4244e+06, 6.4245e+06, 6.4245e+06, 6.4246e+06, 
    6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 6.4249e+06, 6.4249e+06, 
    6.425e+06, 6.4251e+06, 6.4251e+06, 6.4252e+06, 6.4252e+06, 6.4253e+06, 
    6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4256e+06, 6.4256e+06, 6.4257e+06, 
    6.4257e+06, 6.4258e+06, 6.4259e+06, 6.4259e+06, 6.426e+06, 6.426e+06, 
    6.4261e+06, 6.4262e+06, 6.4262e+06, 6.4263e+06, 6.4263e+06, 6.4264e+06, 
    6.4264e+06, 6.4265e+06, 6.4266e+06, 6.4266e+06, 6.4267e+06, 6.4267e+06, 
    6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 6.427e+06, 6.4271e+06, 
    6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 6.4273e+06, 6.4274e+06, 
    6.4275e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 6.4277e+06, 6.4277e+06, 
    6.4278e+06, 6.4279e+06, 6.4279e+06, 6.428e+06, 6.428e+06, 6.4281e+06, 
    6.4282e+06, 6.4282e+06, 6.4283e+06, 6.4284e+06, 6.4284e+06, 6.4285e+06, 
    6.4285e+06, 6.4286e+06, 6.4287e+06, 6.4287e+06, 6.4288e+06, 6.4289e+06, 
    6.4289e+06, 6.429e+06, 6.429e+06, 6.4291e+06, 6.4292e+06, 6.4292e+06, 
    6.4293e+06, 6.4293e+06, 6.4294e+06, 6.4294e+06, 6.4295e+06, 6.4295e+06, 
    6.4296e+06, 6.4297e+06, 6.4297e+06, 6.4298e+06, 6.4298e+06, 6.4299e+06, 
    6.4299e+06, 6.43e+06, 6.4301e+06, 6.4301e+06, 6.4302e+06, 6.4302e+06, 
    6.4303e+06, 6.4304e+06, 6.4304e+06, 6.4305e+06, 6.4305e+06, 6.4306e+06, 
    6.4307e+06, 6.4307e+06, 6.4308e+06, 6.4308e+06, 6.4309e+06, 6.431e+06, 
    6.431e+06, 6.4311e+06, 6.4311e+06, 6.4312e+06, 6.4313e+06, 6.4313e+06, 
    6.4314e+06, 6.4314e+06, 6.4315e+06, 6.4315e+06, 6.4316e+06, 6.4317e+06, 
    6.4317e+06, 6.4318e+06, 6.4318e+06, 6.4319e+06, 6.4319e+06, 6.432e+06, 
    6.432e+06, 6.4321e+06, 6.4321e+06, 6.4322e+06, 6.4322e+06, 6.4323e+06, 
    6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 6.4326e+06, 6.4326e+06, 
    6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4329e+06, 6.4329e+06, 6.433e+06, 
    6.433e+06, 6.4331e+06, 6.4332e+06, 6.4332e+06, 6.4333e+06, 6.4333e+06, 
    6.4334e+06, 6.4335e+06, 6.4335e+06, 6.4336e+06, 6.4336e+06, 6.4337e+06, 
    6.4338e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 6.434e+06, 6.4341e+06, 
    6.4341e+06, 6.4342e+06, 6.4342e+06, 6.4343e+06, 6.4343e+06, 6.4344e+06, 
    6.4344e+06, 6.4345e+06, 6.4346e+06, 6.4346e+06, 6.4347e+06, 6.4347e+06, 
    6.4348e+06, 6.4349e+06, 6.4349e+06, 6.435e+06, 6.435e+06, 6.4351e+06, 
    6.4352e+06, 6.4352e+06, 6.4353e+06, 6.4353e+06, 6.4354e+06, 6.4355e+06, 
    6.4355e+06, 6.4356e+06, 6.4357e+06, 6.4357e+06, 6.4358e+06, 6.4358e+06, 
    6.4359e+06, 6.436e+06, 6.436e+06, 6.4361e+06, 6.4362e+06, 6.4362e+06, 
    6.4363e+06, 6.4364e+06, 6.4364e+06, 6.4365e+06, 6.4366e+06, 6.4366e+06, 
    6.4367e+06, 6.4367e+06, 6.4368e+06, 6.4369e+06, 6.4369e+06, 6.437e+06, 
    6.437e+06, 6.4371e+06, 6.4371e+06, 6.4372e+06, 6.4372e+06, 6.4373e+06, 
    6.4373e+06, 6.4374e+06, 6.4374e+06, 6.4375e+06, 6.4375e+06, 6.4376e+06, 
    6.4376e+06, 6.4377e+06, 6.4377e+06, 6.4378e+06, 6.4379e+06, 6.4379e+06, 
    6.438e+06, 6.438e+06, 6.4381e+06, 6.4381e+06, 6.4382e+06, 6.4382e+06, 
    6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4385e+06, 6.4385e+06, 6.4386e+06, 
    6.4386e+06, 6.4387e+06, 6.4388e+06, 6.4388e+06, 6.4389e+06, 6.439e+06, 
    6.439e+06, 6.4391e+06, 6.4391e+06, 6.4392e+06, 6.4393e+06, 6.4393e+06, 
    6.4394e+06, 6.4395e+06, 6.4395e+06, 6.4396e+06, 6.4396e+06, 6.4397e+06, 
    6.4397e+06, 6.4398e+06, 6.4399e+06, 6.4399e+06, 6.44e+06, 6.44e+06, 
    6.4401e+06, 6.4401e+06, 6.4402e+06, 6.4402e+06, 6.4403e+06, 6.4403e+06, 
    6.4404e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 6.4406e+06, 6.4406e+06, 
    6.4407e+06, 6.4408e+06, 6.4408e+06, 6.4409e+06, 6.4409e+06, 6.441e+06, 
    6.441e+06, 6.4411e+06, 6.4412e+06, 6.4412e+06, 6.4413e+06, 6.4413e+06, 
    6.4414e+06, 6.4415e+06, 6.4415e+06, 6.4416e+06, 6.4417e+06, 6.4417e+06, 
    6.4418e+06, 6.4418e+06, 6.4419e+06, 6.442e+06, 6.442e+06, 6.4421e+06, 
    6.4422e+06, 6.4422e+06, 6.4423e+06, 6.4423e+06, 6.4424e+06, 6.4425e+06, 
    6.4425e+06, 6.4426e+06, 6.4426e+06, 6.4427e+06, 6.4428e+06, 6.4428e+06, 
    6.4429e+06, 6.4429e+06, 6.443e+06, 6.4431e+06, 6.4431e+06, 6.4432e+06, 
    6.4432e+06, 6.4433e+06, 6.4434e+06, 6.4434e+06, 6.4435e+06, 6.4435e+06, 
    6.4436e+06, 6.4437e+06, 6.4437e+06, 6.4438e+06, 6.4438e+06, 6.4439e+06, 
    6.4439e+06, 6.444e+06, 6.444e+06, 6.4441e+06, 6.4441e+06, 6.4442e+06, 
    6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 6.4444e+06, 6.4445e+06, 
    6.4445e+06, 6.4446e+06, 6.4447e+06, 6.4447e+06, 6.4448e+06, 6.4448e+06, 
    6.4449e+06, 6.4449e+06, 6.445e+06, 6.4451e+06, 6.4451e+06, 6.4452e+06, 
    6.4453e+06, 6.4453e+06, 6.4454e+06, 6.4455e+06, 6.4455e+06, 6.4456e+06, 
    6.4456e+06, 6.4457e+06, 6.4458e+06, 6.4458e+06, 6.4459e+06, 6.4459e+06, 
    6.446e+06, 6.4461e+06, 6.4461e+06, 6.4462e+06, 6.4462e+06, 6.4463e+06, 
    6.4463e+06, 6.4464e+06, 6.4464e+06, 6.4465e+06, 6.4465e+06, 6.4466e+06, 
    6.4466e+06, 6.4467e+06, 6.4468e+06, 6.4468e+06, 6.4469e+06, 6.4469e+06, 
    6.447e+06, 6.447e+06, 6.4471e+06, 6.4472e+06, 6.4472e+06, 6.4473e+06, 
    6.4473e+06, 6.4474e+06, 6.4475e+06, 6.4475e+06, 6.4476e+06, 6.4476e+06, 
    6.4477e+06, 6.4478e+06, 6.4478e+06, 6.4479e+06, 6.4479e+06, 6.448e+06, 
    6.4481e+06, 6.4481e+06, 6.4482e+06, 6.4482e+06, 6.4483e+06, 6.4483e+06, 
    6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4486e+06, 6.4486e+06, 6.4487e+06, 
    6.4487e+06, 6.4488e+06, 6.4488e+06, 6.4489e+06, 6.449e+06, 6.449e+06, 
    6.4491e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 6.4493e+06, 6.4494e+06, 
    6.4494e+06, 6.4495e+06, 6.4495e+06, 6.4496e+06, 6.4497e+06, 6.4497e+06, 
    6.4498e+06, 6.4498e+06, 6.4499e+06, 6.45e+06, 6.45e+06, 6.4501e+06, 
    6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 6.4504e+06, 6.4504e+06, 
    6.4505e+06, 6.4505e+06, 6.4506e+06, 6.4507e+06, 6.4507e+06, 6.4508e+06, 
    6.4508e+06, 6.4509e+06, 6.4509e+06, 6.451e+06, 6.4511e+06, 6.4511e+06, 
    6.4512e+06, 6.4512e+06, 6.4513e+06, 6.4514e+06, 6.4514e+06, 6.4515e+06, 
    6.4515e+06, 6.4516e+06, 6.4517e+06, 6.4517e+06, 6.4518e+06, 6.4518e+06, 
    6.4519e+06, 6.452e+06, 6.452e+06, 6.4521e+06, 6.4521e+06, 6.4522e+06, 
    6.4522e+06, 6.4523e+06, 6.4524e+06, 6.4524e+06, 6.4525e+06, 6.4525e+06, 
    6.4526e+06, 6.4526e+06, 6.4527e+06, 6.4527e+06, 6.4528e+06, 6.4529e+06, 
    6.4529e+06, 6.453e+06, 6.453e+06, 6.4531e+06, 6.4531e+06, 6.4532e+06, 
    6.4533e+06, 6.4533e+06, 6.4534e+06, 6.4535e+06, 6.4535e+06, 6.4536e+06, 
    6.4536e+06, 6.4537e+06, 6.4538e+06, 6.4538e+06, 6.4539e+06, 6.4539e+06, 
    6.454e+06, 6.454e+06, 6.4541e+06, 6.4541e+06, 6.4542e+06, 6.4543e+06, 
    6.4543e+06, 6.4544e+06, 6.4544e+06, 6.4545e+06, 6.4545e+06, 6.4546e+06, 
    6.4546e+06, 6.4547e+06, 6.4547e+06, 6.4548e+06, 6.4548e+06, 6.4549e+06, 
    6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 6.4551e+06, 6.4552e+06, 
    6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 6.4555e+06, 6.4556e+06, 
    6.4556e+06, 6.4557e+06, 6.4558e+06, 6.4558e+06, 6.4559e+06, 6.456e+06, 
    6.456e+06, 6.4561e+06, 6.4561e+06, 6.4562e+06, 6.4563e+06, 6.4563e+06, 
    6.4564e+06, 6.4564e+06, 6.4565e+06, 6.4566e+06, 6.4566e+06, 6.4567e+06, 
    6.4567e+06, 6.4568e+06, 6.4568e+06, 6.4569e+06, 6.4569e+06,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 6.3923e+06, 6.3923e+06, 
    6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 6.3924e+06, 6.3924e+06, 
    6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 6.3926e+06, 6.3926e+06, 
    6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 6.3927e+06, 
    6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 
    6.3929e+06, 6.393e+06, 6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 
    6.3931e+06, 6.3931e+06, 6.3932e+06, 6.3932e+06, 6.3932e+06, 6.3933e+06, 
    6.3933e+06, 6.3933e+06, 6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 
    6.3935e+06, 6.3935e+06, 6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 
    6.3937e+06, 6.3937e+06, 6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 
    6.3938e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 6.3939e+06, 
    6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.3941e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 6.3944e+06, 
    6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 6.3946e+06, 
    6.3947e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 6.3949e+06, 
    6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 6.3951e+06, 6.3951e+06, 
    6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3953e+06, 6.3953e+06, 6.3953e+06, 
    6.3954e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 6.3955e+06, 6.3956e+06, 
    6.3956e+06, 6.3956e+06, 6.3957e+06, 6.3957e+06, 6.3957e+06, 6.3958e+06, 
    6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 6.396e+06, 6.396e+06, 
    6.396e+06, 6.3961e+06, 6.3961e+06, 6.3961e+06, 6.3962e+06, 6.3962e+06, 
    6.3963e+06, 6.3963e+06, 6.3963e+06, 6.3964e+06, 6.3964e+06, 6.3964e+06, 
    6.3965e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 6.3966e+06, 6.3966e+06, 
    6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 6.3968e+06, 6.3969e+06, 
    6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 6.397e+06, 6.3971e+06, 
    6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 6.3973e+06, 6.3973e+06, 
    6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3975e+06, 6.3975e+06, 6.3975e+06, 
    6.3976e+06, 6.3976e+06, 6.3977e+06, 6.3977e+06, 6.3977e+06, 6.3978e+06, 
    6.3978e+06, 6.3979e+06, 6.3979e+06, 6.398e+06, 6.398e+06, 6.3981e+06, 
    6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 6.3983e+06, 6.3983e+06, 
    6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 6.3986e+06, 6.3986e+06, 
    6.3987e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 6.3988e+06, 6.3989e+06, 
    6.3989e+06, 6.399e+06, 6.399e+06, 6.399e+06, 6.3991e+06, 6.3991e+06, 
    6.3992e+06, 6.3992e+06, 6.3992e+06, 6.3993e+06, 6.3993e+06, 6.3994e+06, 
    6.3994e+06, 6.3994e+06, 6.3995e+06, 6.3995e+06, 6.3995e+06, 6.3996e+06, 
    6.3996e+06, 6.3997e+06, 6.3997e+06, 6.3997e+06, 6.3998e+06, 6.3998e+06, 
    6.3999e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 6.4e+06, 6.4001e+06, 
    6.4001e+06, 6.4002e+06, 6.4002e+06, 6.4003e+06, 6.4003e+06, 6.4004e+06, 
    6.4004e+06, 6.4005e+06, 6.4005e+06, 6.4005e+06, 6.4006e+06, 6.4006e+06, 
    6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 6.4009e+06, 6.4009e+06, 
    6.401e+06, 6.401e+06, 6.4011e+06, 6.4011e+06, 6.4011e+06, 6.4012e+06, 
    6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4014e+06, 6.4014e+06, 6.4015e+06, 
    6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 6.4017e+06, 6.4017e+06, 
    6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 6.402e+06, 6.402e+06, 
    6.4021e+06, 6.4021e+06, 6.4022e+06, 6.4022e+06, 6.4023e+06, 6.4023e+06, 
    6.4024e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 6.4026e+06, 6.4026e+06, 
    6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 6.4029e+06, 6.4029e+06, 
    6.403e+06, 6.403e+06, 6.4031e+06, 6.4031e+06, 6.4032e+06, 6.4032e+06, 
    6.4033e+06, 6.4033e+06, 6.4034e+06, 6.4034e+06, 6.4035e+06, 6.4035e+06, 
    6.4036e+06, 6.4036e+06, 6.4037e+06, 6.4037e+06, 6.4038e+06, 6.4038e+06, 
    6.4039e+06, 6.4039e+06, 6.404e+06, 6.404e+06, 6.4041e+06, 6.4041e+06, 
    6.4042e+06, 6.4042e+06, 6.4043e+06, 6.4043e+06, 6.4044e+06, 6.4044e+06, 
    6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 6.4047e+06, 6.4048e+06, 
    6.4048e+06, 6.4049e+06, 6.4049e+06, 6.405e+06, 6.405e+06, 6.4051e+06, 
    6.4051e+06, 6.4052e+06, 6.4052e+06, 6.4053e+06, 6.4054e+06, 6.4054e+06, 
    6.4055e+06, 6.4055e+06, 6.4056e+06, 6.4056e+06, 6.4057e+06, 6.4057e+06, 
    6.4058e+06, 6.4058e+06, 6.4059e+06, 6.406e+06, 6.406e+06, 6.4061e+06, 
    6.4061e+06, 6.4062e+06, 6.4062e+06, 6.4063e+06, 6.4063e+06, 6.4064e+06, 
    6.4064e+06, 6.4065e+06, 6.4065e+06, 6.4065e+06, 6.4066e+06, 6.4066e+06, 
    6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 6.4069e+06, 6.4069e+06, 
    6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 6.4072e+06, 6.4072e+06, 
    6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 6.4075e+06, 6.4076e+06, 
    6.4076e+06, 6.4077e+06, 6.4077e+06, 6.4078e+06, 6.4078e+06, 6.4079e+06, 
    6.408e+06, 6.408e+06, 6.4081e+06, 6.4081e+06, 6.4082e+06, 6.4082e+06, 
    6.4083e+06, 6.4084e+06, 6.4084e+06, 6.4085e+06, 6.4085e+06, 6.4086e+06, 
    6.4086e+06, 6.4087e+06, 6.4087e+06, 6.4088e+06, 6.4088e+06, 6.4089e+06, 
    6.409e+06, 6.409e+06, 6.4091e+06, 6.4091e+06, 6.4092e+06, 6.4092e+06, 
    6.4093e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 6.4095e+06, 6.4096e+06, 
    6.4096e+06, 6.4097e+06, 6.4097e+06, 6.4098e+06, 6.4098e+06, 6.4099e+06, 
    6.41e+06, 6.41e+06, 6.4101e+06, 6.4101e+06, 6.4102e+06, 6.4102e+06, 
    6.4103e+06, 6.4104e+06, 6.4104e+06, 6.4105e+06, 6.4105e+06, 6.4106e+06, 
    6.4106e+06, 6.4107e+06, 6.4107e+06, 6.4108e+06, 6.4108e+06, 6.4109e+06, 
    6.411e+06, 6.411e+06, 6.4111e+06, 6.4111e+06, 6.4112e+06, 6.4112e+06, 
    6.4113e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 6.4115e+06, 6.4115e+06, 
    6.4116e+06, 6.4117e+06, 6.4117e+06, 6.4118e+06, 6.4118e+06, 6.4119e+06, 
    6.4119e+06, 6.412e+06, 6.4121e+06, 6.4121e+06, 6.4122e+06, 6.4122e+06, 
    6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4125e+06, 6.4125e+06, 6.4126e+06, 
    6.4126e+06, 6.4127e+06, 6.4127e+06, 6.4128e+06, 6.4129e+06, 6.4129e+06, 
    6.413e+06, 6.413e+06, 6.4131e+06, 6.4131e+06, 6.4132e+06, 6.4132e+06, 
    6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 6.4135e+06, 6.4136e+06, 
    6.4136e+06, 6.4137e+06, 6.4137e+06, 6.4138e+06, 6.4138e+06, 6.4139e+06, 
    6.4139e+06, 6.414e+06, 6.4141e+06, 6.4141e+06, 6.4142e+06, 6.4142e+06, 
    6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4145e+06, 6.4145e+06, 6.4146e+06, 
    6.4146e+06, 6.4147e+06, 6.4148e+06, 6.4148e+06, 6.4149e+06, 6.4149e+06, 
    6.415e+06, 6.4151e+06, 6.4151e+06, 6.4152e+06, 6.4152e+06, 6.4153e+06, 
    6.4154e+06, 6.4154e+06, 6.4155e+06, 6.4156e+06, 6.4156e+06, 6.4157e+06, 
    6.4157e+06, 6.4158e+06, 6.4158e+06, 6.4159e+06, 6.416e+06, 6.416e+06, 
    6.4161e+06, 6.4161e+06, 6.4162e+06, 6.4162e+06, 6.4163e+06, 6.4164e+06, 
    6.4164e+06, 6.4165e+06, 6.4165e+06, 6.4166e+06, 6.4166e+06, 6.4167e+06, 
    6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 6.4169e+06, 6.417e+06, 
    6.4171e+06, 6.4171e+06, 6.4172e+06, 6.4172e+06, 6.4173e+06, 6.4173e+06, 
    6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 6.4176e+06, 6.4177e+06, 
    6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 6.4179e+06, 6.418e+06, 
    6.4181e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 6.4183e+06, 6.4183e+06, 
    6.4184e+06, 6.4185e+06, 6.4185e+06, 6.4186e+06, 6.4186e+06, 6.4187e+06, 
    6.4187e+06, 6.4188e+06, 6.4189e+06, 6.4189e+06, 6.419e+06, 6.419e+06, 
    6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4193e+06, 6.4193e+06, 6.4194e+06, 
    6.4194e+06, 6.4195e+06, 6.4196e+06, 6.4196e+06, 6.4197e+06, 6.4197e+06, 
    6.4198e+06, 6.4199e+06, 6.4199e+06, 6.42e+06, 6.42e+06, 6.4201e+06, 
    6.4202e+06, 6.4202e+06, 6.4203e+06, 6.4203e+06, 6.4204e+06, 6.4205e+06, 
    6.4205e+06, 6.4206e+06, 6.4206e+06, 6.4207e+06, 6.4207e+06, 6.4208e+06, 
    6.4209e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 6.4211e+06, 6.4212e+06, 
    6.4212e+06, 6.4213e+06, 6.4213e+06, 6.4214e+06, 6.4214e+06, 6.4215e+06, 
    6.4216e+06, 6.4216e+06, 6.4217e+06, 6.4217e+06, 6.4218e+06, 6.4219e+06, 
    6.4219e+06, 6.422e+06, 6.422e+06, 6.4221e+06, 6.4222e+06, 6.4222e+06, 
    6.4223e+06, 6.4224e+06, 6.4224e+06, 6.4225e+06, 6.4226e+06, 6.4226e+06, 
    6.4227e+06, 6.4228e+06, 6.4228e+06, 6.4229e+06, 6.4229e+06, 6.423e+06, 
    6.4231e+06, 6.4231e+06, 6.4232e+06, 6.4232e+06, 6.4233e+06, 6.4234e+06, 
    6.4234e+06, 6.4235e+06, 6.4235e+06, 6.4236e+06, 6.4236e+06, 6.4237e+06, 
    6.4237e+06, 6.4238e+06, 6.4238e+06, 6.4239e+06, 6.4239e+06, 6.424e+06, 
    6.424e+06, 6.4241e+06, 6.4241e+06, 6.4242e+06, 6.4242e+06, 6.4243e+06, 
    6.4243e+06, 6.4244e+06, 6.4244e+06, 6.4245e+06, 6.4245e+06, 6.4246e+06, 
    6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 6.4249e+06, 6.4249e+06, 
    6.425e+06, 6.4251e+06, 6.4251e+06, 6.4252e+06, 6.4252e+06, 6.4253e+06, 
    6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4256e+06, 6.4256e+06, 6.4257e+06, 
    6.4257e+06, 6.4258e+06, 6.4259e+06, 6.4259e+06, 6.426e+06, 6.426e+06, 
    6.4261e+06, 6.4262e+06, 6.4262e+06, 6.4263e+06, 6.4263e+06, 6.4264e+06, 
    6.4264e+06, 6.4265e+06, 6.4266e+06, 6.4266e+06, 6.4267e+06, 6.4267e+06, 
    6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 6.427e+06, 6.4271e+06, 
    6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 6.4273e+06, 6.4274e+06, 
    6.4275e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 6.4277e+06, 6.4277e+06, 
    6.4278e+06, 6.4279e+06, 6.4279e+06, 6.428e+06, 6.428e+06, 6.4281e+06, 
    6.4282e+06, 6.4282e+06, 6.4283e+06, 6.4284e+06, 6.4284e+06, 6.4285e+06, 
    6.4285e+06, 6.4286e+06, 6.4287e+06, 6.4287e+06, 6.4288e+06, 6.4289e+06, 
    6.4289e+06, 6.429e+06, 6.429e+06, 6.4291e+06, 6.4292e+06, 6.4292e+06, 
    6.4293e+06, 6.4293e+06, 6.4294e+06, 6.4294e+06, 6.4295e+06, 6.4295e+06, 
    6.4296e+06, 6.4297e+06, 6.4297e+06, 6.4298e+06, 6.4298e+06, 6.4299e+06, 
    6.4299e+06, 6.43e+06, 6.4301e+06, 6.4301e+06, 6.4302e+06, 6.4302e+06, 
    6.4303e+06, 6.4304e+06, 6.4304e+06, 6.4305e+06, 6.4305e+06, 6.4306e+06, 
    6.4307e+06, 6.4307e+06, 6.4308e+06, 6.4308e+06, 6.4309e+06, 6.431e+06, 
    6.431e+06, 6.4311e+06, 6.4311e+06, 6.4312e+06, 6.4313e+06, 6.4313e+06, 
    6.4314e+06, 6.4314e+06, 6.4315e+06, 6.4315e+06, 6.4316e+06, 6.4317e+06, 
    6.4317e+06, 6.4318e+06, 6.4318e+06, 6.4319e+06, 6.4319e+06, 6.432e+06, 
    6.432e+06, 6.4321e+06, 6.4321e+06, 6.4322e+06, 6.4322e+06, 6.4323e+06, 
    6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 6.4326e+06, 6.4326e+06, 
    6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4329e+06, 6.4329e+06, 6.433e+06, 
    6.433e+06, 6.4331e+06, 6.4332e+06, 6.4332e+06, 6.4333e+06, 6.4333e+06, 
    6.4334e+06, 6.4335e+06, 6.4335e+06, 6.4336e+06, 6.4336e+06, 6.4337e+06, 
    6.4338e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 6.434e+06, 6.4341e+06, 
    6.4341e+06, 6.4342e+06, 6.4342e+06, 6.4343e+06, 6.4343e+06, 6.4344e+06, 
    6.4344e+06, 6.4345e+06, 6.4346e+06, 6.4346e+06, 6.4347e+06, 6.4347e+06, 
    6.4348e+06, 6.4349e+06, 6.4349e+06, 6.435e+06, 6.435e+06, 6.4351e+06, 
    6.4352e+06, 6.4352e+06, 6.4353e+06, 6.4353e+06, 6.4354e+06, 6.4355e+06, 
    6.4355e+06, 6.4356e+06, 6.4357e+06, 6.4357e+06, 6.4358e+06, 6.4358e+06, 
    6.4359e+06, 6.436e+06, 6.436e+06, 6.4361e+06, 6.4362e+06, 6.4362e+06, 
    6.4363e+06, 6.4364e+06, 6.4364e+06, 6.4365e+06, 6.4366e+06, 6.4366e+06, 
    6.4367e+06, 6.4367e+06, 6.4368e+06, 6.4369e+06, 6.4369e+06, 6.437e+06, 
    6.437e+06, 6.4371e+06, 6.4371e+06, 6.4372e+06, 6.4372e+06, 6.4373e+06, 
    6.4373e+06, 6.4374e+06, 6.4374e+06, 6.4375e+06, 6.4375e+06, 6.4376e+06, 
    6.4376e+06, 6.4377e+06, 6.4377e+06, 6.4378e+06, 6.4379e+06, 6.4379e+06, 
    6.438e+06, 6.438e+06, 6.4381e+06, 6.4381e+06, 6.4382e+06, 6.4382e+06, 
    6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4385e+06, 6.4385e+06, 6.4386e+06, 
    6.4386e+06, 6.4387e+06, 6.4388e+06, 6.4388e+06, 6.4389e+06, 6.439e+06, 
    6.439e+06, 6.4391e+06, 6.4391e+06, 6.4392e+06, 6.4393e+06, 6.4393e+06, 
    6.4394e+06, 6.4395e+06, 6.4395e+06, 6.4396e+06, 6.4396e+06, 6.4397e+06, 
    6.4397e+06, 6.4398e+06, 6.4399e+06, 6.4399e+06, 6.44e+06, 6.44e+06, 
    6.4401e+06, 6.4401e+06, 6.4402e+06, 6.4402e+06, 6.4403e+06, 6.4403e+06, 
    6.4404e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 6.4406e+06, 6.4406e+06, 
    6.4407e+06, 6.4408e+06, 6.4408e+06, 6.4409e+06, 6.4409e+06, 6.441e+06, 
    6.441e+06, 6.4411e+06, 6.4412e+06, 6.4412e+06, 6.4413e+06, 6.4413e+06, 
    6.4414e+06, 6.4415e+06, 6.4415e+06, 6.4416e+06, 6.4417e+06, 6.4417e+06, 
    6.4418e+06, 6.4418e+06, 6.4419e+06, 6.442e+06, 6.442e+06, 6.4421e+06, 
    6.4422e+06, 6.4422e+06, 6.4423e+06, 6.4423e+06, 6.4424e+06, 6.4425e+06, 
    6.4425e+06, 6.4426e+06, 6.4426e+06, 6.4427e+06, 6.4428e+06, 6.4428e+06, 
    6.4429e+06, 6.4429e+06, 6.443e+06, 6.4431e+06, 6.4431e+06, 6.4432e+06, 
    6.4432e+06, 6.4433e+06, 6.4434e+06, 6.4434e+06, 6.4435e+06, 6.4435e+06, 
    6.4436e+06, 6.4437e+06, 6.4437e+06, 6.4438e+06, 6.4438e+06, 6.4439e+06, 
    6.4439e+06, 6.444e+06, 6.444e+06, 6.4441e+06, 6.4441e+06, 6.4442e+06, 
    6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 6.4444e+06, 6.4445e+06, 
    6.4445e+06, 6.4446e+06, 6.4447e+06, 6.4447e+06, 6.4448e+06, 6.4448e+06, 
    6.4449e+06, 6.4449e+06, 6.445e+06, 6.4451e+06, 6.4451e+06, 6.4452e+06, 
    6.4453e+06, 6.4453e+06, 6.4454e+06, 6.4455e+06, 6.4455e+06, 6.4456e+06, 
    6.4456e+06, 6.4457e+06, 6.4458e+06, 6.4458e+06, 6.4459e+06, 6.4459e+06, 
    6.446e+06, 6.4461e+06, 6.4461e+06, 6.4462e+06, 6.4462e+06, 6.4463e+06, 
    6.4463e+06, 6.4464e+06, 6.4464e+06, 6.4465e+06, 6.4465e+06, 6.4466e+06, 
    6.4466e+06, 6.4467e+06, 6.4468e+06, 6.4468e+06, 6.4469e+06, 6.4469e+06, 
    6.447e+06, 6.447e+06, 6.4471e+06, 6.4472e+06, 6.4472e+06, 6.4473e+06, 
    6.4473e+06, 6.4474e+06, 6.4475e+06, 6.4475e+06, 6.4476e+06, 6.4476e+06, 
    6.4477e+06, 6.4478e+06, 6.4478e+06, 6.4479e+06, 6.4479e+06, 6.448e+06, 
    6.4481e+06, 6.4481e+06, 6.4482e+06, 6.4482e+06, 6.4483e+06, 6.4483e+06, 
    6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4486e+06, 6.4486e+06, 6.4487e+06, 
    6.4487e+06, 6.4488e+06, 6.4488e+06, 6.4489e+06, 6.449e+06, 6.449e+06, 
    6.4491e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 6.4493e+06, 6.4494e+06, 
    6.4494e+06, 6.4495e+06, 6.4495e+06, 6.4496e+06, 6.4497e+06, 6.4497e+06, 
    6.4498e+06, 6.4498e+06, 6.4499e+06, 6.45e+06, 6.45e+06, 6.4501e+06, 
    6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 6.4504e+06, 6.4504e+06, 
    6.4505e+06, 6.4505e+06, 6.4506e+06, 6.4507e+06, 6.4507e+06, 6.4508e+06, 
    6.4508e+06, 6.4509e+06, 6.4509e+06, 6.451e+06, 6.4511e+06, 6.4511e+06, 
    6.4512e+06, 6.4512e+06, 6.4513e+06, 6.4514e+06, 6.4514e+06, 6.4515e+06, 
    6.4515e+06, 6.4516e+06, 6.4517e+06, 6.4517e+06, 6.4518e+06, 6.4518e+06, 
    6.4519e+06, 6.452e+06, 6.452e+06, 6.4521e+06, 6.4521e+06, 6.4522e+06, 
    6.4522e+06, 6.4523e+06, 6.4524e+06, 6.4524e+06, 6.4525e+06, 6.4525e+06, 
    6.4526e+06, 6.4526e+06, 6.4527e+06, 6.4527e+06, 6.4528e+06, 6.4529e+06, 
    6.4529e+06, 6.453e+06, 6.453e+06, 6.4531e+06, 6.4531e+06, 6.4532e+06, 
    6.4533e+06, 6.4533e+06, 6.4534e+06, 6.4535e+06, 6.4535e+06, 6.4536e+06, 
    6.4536e+06, 6.4537e+06, 6.4538e+06, 6.4538e+06, 6.4539e+06, 6.4539e+06, 
    6.454e+06, 6.454e+06, 6.4541e+06, 6.4541e+06, 6.4542e+06, 6.4543e+06, 
    6.4543e+06, 6.4544e+06, 6.4544e+06, 6.4545e+06, 6.4545e+06, 6.4546e+06, 
    6.4546e+06, 6.4547e+06, 6.4547e+06, 6.4548e+06, 6.4548e+06, 6.4549e+06, 
    6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 6.4551e+06, 6.4552e+06, 
    6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 6.4555e+06, 6.4556e+06, 
    6.4556e+06, 6.4557e+06, 6.4558e+06, 6.4558e+06, 6.4559e+06, 6.456e+06, 
    6.456e+06, 6.4561e+06, 6.4561e+06, 6.4562e+06, 6.4563e+06, 6.4563e+06, 
    6.4564e+06, 6.4564e+06, 6.4565e+06, 6.4566e+06, 6.4566e+06, 6.4567e+06, 
    6.4567e+06, 6.4568e+06, 6.4568e+06, 6.4569e+06, 6.4569e+06 ;

 impact =
  6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.377e+06, 6.377e+06, 
    6.377e+06, 6.377e+06, 6.3771e+06, 6.3771e+06, 6.3772e+06, 6.3772e+06, 
    6.3772e+06, 6.3773e+06, 6.3773e+06, 6.3774e+06, 6.3774e+06, 6.3775e+06, 
    6.3775e+06, 6.3775e+06, 6.3776e+06, 6.3776e+06, 6.3777e+06, 6.3777e+06, 
    6.3777e+06, 6.3777e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3782e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 
    6.3784e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3786e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.3789e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3786e+06, 6.3786e+06, 6.3786e+06, 
    6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3784e+06, 
    6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 
    6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3782e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3781e+06, 6.3781e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 6.3784e+06, 
    6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3796e+06, 
    6.3796e+06, 6.3796e+06, 6.3797e+06, 6.3797e+06, 6.3798e+06, 6.3798e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.38e+06, 
    6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3798e+06, 6.3798e+06, 
    6.3798e+06, 6.3798e+06, 6.3797e+06, 6.3797e+06, 6.3796e+06, 6.3796e+06, 
    6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3794e+06, 6.3794e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3805e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3805e+06, 6.3805e+06, 
    6.3805e+06, 6.3805e+06, 6.3805e+06, 6.3806e+06, 6.3806e+06, 6.3806e+06, 
    6.3807e+06, 6.3807e+06, 6.3807e+06, 6.3808e+06, 6.3808e+06, 6.3808e+06, 
    6.3809e+06, 6.3809e+06, 6.3809e+06, 6.381e+06, 6.381e+06, 6.381e+06, 
    6.381e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 
    6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 
    6.3815e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 
    6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 
    6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 
    6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 
    6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 
    6.382e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 
    6.3821e+06, 6.3821e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 
    6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3823e+06, 6.3823e+06, 
    6.3823e+06, 6.3823e+06, 6.3823e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 
    6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3825e+06, 6.3825e+06, 
    6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 
    6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3827e+06, 
    6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3828e+06, 6.3828e+06, 
    6.3828e+06, 6.3828e+06, 6.3828e+06, 6.3829e+06, 6.3829e+06, 6.3829e+06, 
    6.3829e+06, 6.3829e+06, 6.383e+06, 6.383e+06, 6.383e+06, 6.383e+06, 
    6.383e+06, 6.383e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 
    6.3831e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 
    6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 
    6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3837e+06, 
    6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3838e+06, 
    6.3838e+06, 6.3838e+06, 6.3838e+06, 6.3839e+06, 6.3839e+06, 6.3839e+06, 
    6.3839e+06, 6.3839e+06, 6.3839e+06, 6.384e+06, 6.384e+06, 6.384e+06, 
    6.384e+06, 6.384e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 
    6.3841e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3843e+06, 
    6.3843e+06, 6.3843e+06, 6.3843e+06, 6.3844e+06, 6.3844e+06, 6.3844e+06, 
    6.3844e+06, 6.3845e+06, 6.3845e+06, 6.3845e+06, 6.3846e+06, 6.3846e+06, 
    6.3846e+06, 6.3846e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 
    6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3849e+06, 
    6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.385e+06, 
    6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 
    6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 
    6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3853e+06, 
    6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3854e+06, 
    6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3855e+06, 6.3855e+06, 
    6.3855e+06, 6.3855e+06, 6.3855e+06, 6.3856e+06, 6.3856e+06, 6.3856e+06, 
    6.3856e+06, 6.3856e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 
    6.3857e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3859e+06, 
    6.3859e+06, 6.3859e+06, 6.3859e+06, 6.3859e+06, 6.386e+06, 6.386e+06, 
    6.386e+06, 6.386e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.3951e+06, 6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3962e+06, 6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 
    6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3975e+06, 6.3975e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 
    6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 
    6.3983e+06, 6.3983e+06, 6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3986e+06, 6.3986e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3993e+06, 6.3993e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3995e+06, 
    6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 
    6.4006e+06, 6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 
    6.4008e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 
    6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 
    6.4017e+06, 6.4017e+06, 6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 
    6.4029e+06, 6.4029e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4037e+06, 
    6.4037e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 
    6.404e+06, 6.4041e+06, 6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 
    6.405e+06, 6.405e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 
    6.406e+06, 6.406e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 
    6.4063e+06, 6.4063e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 6.4065e+06, 
    6.4066e+06, 6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 
    6.4069e+06, 6.4069e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4072e+06, 6.4072e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4079e+06, 6.4079e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4082e+06, 6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 6.4084e+06, 
    6.4085e+06, 6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4088e+06, 
    6.4088e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.4091e+06, 
    6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4095e+06, 6.4095e+06, 6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 
    6.4098e+06, 6.4099e+06, 6.4099e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 
    6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4107e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 6.411e+06, 6.4111e+06, 
    6.4111e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 
    6.4115e+06, 6.4115e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4119e+06, 6.4119e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 
    6.4121e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4124e+06, 
    6.4125e+06, 6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4128e+06, 
    6.4128e+06, 6.4129e+06, 6.4129e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 6.4138e+06, 
    6.4138e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.4141e+06, 
    6.4141e+06, 6.4142e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 
    6.4148e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.4151e+06, 6.4151e+06, 
    6.4152e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4155e+06, 
    6.4156e+06, 6.4156e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4159e+06, 
    6.4159e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 6.4161e+06, 6.4162e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 6.4165e+06, 
    6.4166e+06, 6.4166e+06, 6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 6.4172e+06, 
    6.4172e+06, 6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 
    6.4179e+06, 6.418e+06, 6.418e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 
    6.4183e+06, 6.4183e+06, 6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 6.4189e+06, 
    6.419e+06, 6.419e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 6.42e+06, 
    6.42e+06, 6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 
    6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 6.4206e+06, 6.4207e+06, 
    6.4207e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 
    6.4211e+06, 6.4211e+06, 6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 6.4217e+06, 
    6.4218e+06, 6.4218e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.4221e+06, 
    6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 6.4227e+06, 6.4228e+06, 
    6.4229e+06, 6.4229e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 6.4232e+06, 
    6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 6.4238e+06, 
    6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 6.4241e+06, 6.4241e+06, 
    6.4242e+06, 6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4245e+06, 
    6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 6.4252e+06, 
    6.4252e+06, 6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4258e+06, 6.4258e+06, 6.4259e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 6.4262e+06, 
    6.4263e+06, 6.4264e+06, 6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 
    6.4266e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 
    6.427e+06, 6.427e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 
    6.4277e+06, 6.4277e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 6.4283e+06, 6.4283e+06, 
    6.4284e+06, 6.4284e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4287e+06, 
    6.4288e+06, 6.4288e+06, 6.4289e+06, 6.4289e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 6.4294e+06, 
    6.4295e+06, 6.4295e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.43e+06, 6.43e+06, 6.4301e+06, 
    6.4301e+06, 6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 6.4312e+06, 
    6.4312e+06, 6.4313e+06, 6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4318e+06, 6.4318e+06, 
    6.4319e+06, 6.4319e+06, 6.432e+06, 6.432e+06, 6.4321e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 
    6.4326e+06, 6.4326e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 6.4331e+06, 6.4332e+06, 
    6.4333e+06, 6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4336e+06, 
    6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4343e+06, 
    6.4343e+06, 6.4344e+06, 6.4344e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 6.4349e+06, 
    6.435e+06, 6.4351e+06, 6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 
    6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4356e+06, 6.4357e+06, 
    6.4357e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 6.436e+06, 
    6.4361e+06, 6.4362e+06, 6.4362e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 
    6.4368e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 6.4371e+06, 
    6.4372e+06, 6.4372e+06, 6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 
    6.4375e+06, 6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4378e+06, 
    6.4378e+06, 6.4379e+06, 6.4379e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4384e+06, 
    6.4385e+06, 6.4386e+06, 6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.4391e+06, 6.4392e+06, 
    6.4392e+06, 6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4395e+06, 6.4395e+06, 
    6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 
    6.4399e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4402e+06, 
    6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 
    6.4406e+06, 6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4409e+06, 
    6.4409e+06, 6.441e+06, 6.441e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 6.4416e+06, 
    6.4416e+06, 6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.4421e+06, 6.4421e+06, 6.4422e+06, 6.4422e+06, 6.4423e+06, 
    6.4423e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4427e+06, 6.4428e+06, 6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4433e+06, 6.4434e+06, 
    6.4434e+06, 6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 6.444e+06, 6.444e+06, 
    6.4441e+06, 6.4441e+06, 6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 
    6.4444e+06, 6.4445e+06, 6.4445e+06, 6.4446e+06, 6.4446e+06, 6.4447e+06, 
    6.4447e+06, 6.4448e+06, 6.4449e+06, 6.4449e+06, 6.445e+06, 6.445e+06, 
    6.4451e+06, 6.4452e+06, 6.4452e+06, 6.4453e+06, 6.4453e+06, 6.4454e+06, 
    6.4455e+06, 6.4455e+06, 6.4456e+06, 6.4457e+06, 6.4457e+06, 6.4458e+06, 
    6.4458e+06, 6.4459e+06, 6.4459e+06, 6.446e+06, 6.4461e+06, 6.4461e+06, 
    6.4462e+06, 6.4462e+06, 6.4463e+06, 6.4463e+06, 6.4464e+06, 6.4465e+06, 
    6.4465e+06, 6.4466e+06, 6.4466e+06, 6.4467e+06, 6.4467e+06, 6.4468e+06, 
    6.4468e+06, 6.4469e+06, 6.447e+06, 6.447e+06, 6.4471e+06, 6.4471e+06, 
    6.4472e+06, 6.4472e+06, 6.4473e+06, 6.4474e+06, 6.4474e+06, 6.4475e+06, 
    6.4475e+06, 6.4476e+06, 6.4477e+06, 6.4477e+06, 6.4478e+06, 6.4478e+06, 
    6.4479e+06, 6.448e+06, 6.448e+06, 6.4481e+06, 6.4481e+06, 6.4482e+06, 
    6.4482e+06, 6.4483e+06, 6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4485e+06, 
    6.4486e+06, 6.4486e+06, 6.4487e+06, 6.4487e+06, 6.4488e+06, 6.4489e+06, 
    6.4489e+06, 6.449e+06, 6.449e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 
    6.4493e+06, 6.4493e+06, 6.4494e+06, 6.4494e+06, 6.4495e+06, 6.4496e+06, 
    6.4496e+06, 6.4497e+06, 6.4497e+06, 6.4498e+06, 6.4499e+06, 6.4499e+06, 
    6.45e+06, 6.45e+06, 6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 
    6.4503e+06, 6.4504e+06, 6.4504e+06, 6.4505e+06, 6.4506e+06, 6.4506e+06, 
    6.4507e+06, 6.4507e+06, 6.4508e+06, 6.4508e+06, 6.4509e+06, 6.451e+06, 
    6.451e+06, 6.4511e+06, 6.4511e+06, 6.4512e+06, 6.4513e+06, 6.4513e+06, 
    6.4514e+06, 6.4514e+06, 6.4515e+06, 6.4516e+06, 6.4516e+06, 6.4517e+06, 
    6.4517e+06, 6.4518e+06, 6.4518e+06, 6.4519e+06, 6.452e+06, 6.452e+06, 
    6.4521e+06, 6.4521e+06, 6.4522e+06, 6.4522e+06, 6.4523e+06, 6.4524e+06, 
    6.4524e+06, 6.4525e+06, 6.4525e+06, 6.4526e+06, 6.4526e+06, 6.4527e+06, 
    6.4527e+06, 6.4528e+06, 6.4529e+06, 6.4529e+06, 6.453e+06, 6.453e+06, 
    6.4531e+06, 6.4532e+06, 6.4532e+06, 6.4533e+06, 6.4533e+06, 6.4534e+06, 
    6.4535e+06, 6.4535e+06, 6.4536e+06, 6.4536e+06, 6.4537e+06, 6.4538e+06, 
    6.4538e+06, 6.4539e+06, 6.4539e+06, 6.454e+06, 6.454e+06, 6.4541e+06, 
    6.4541e+06, 6.4542e+06, 6.4543e+06, 6.4543e+06, 6.4544e+06, 6.4544e+06, 
    6.4545e+06, 6.4545e+06, 6.4546e+06, 6.4546e+06, 6.4547e+06, 6.4547e+06, 
    6.4548e+06, 6.4548e+06, 6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 
    6.4551e+06, 6.4552e+06, 6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 
    6.4555e+06, 6.4555e+06, 6.4556e+06, 6.4557e+06, 6.4557e+06, 6.4558e+06, 
    6.4559e+06, 6.4559e+06, 6.456e+06, 6.456e+06, 6.4561e+06, 6.4562e+06, 
    6.4562e+06, 6.4563e+06, 6.4563e+06, 6.4564e+06, 6.4565e+06, 6.4565e+06, 
    6.4566e+06, 6.4566e+06, 6.4567e+06, 6.4567e+06, 6.4568e+06, 6.4568e+06, 
    6.4569e+06,
  6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 6.3768e+06, 
    6.3769e+06, 6.3769e+06, 6.3769e+06, 6.3769e+06, 6.377e+06, 6.377e+06, 
    6.377e+06, 6.377e+06, 6.3771e+06, 6.3771e+06, 6.3772e+06, 6.3772e+06, 
    6.3772e+06, 6.3773e+06, 6.3773e+06, 6.3774e+06, 6.3774e+06, 6.3775e+06, 
    6.3775e+06, 6.3775e+06, 6.3776e+06, 6.3776e+06, 6.3777e+06, 6.3777e+06, 
    6.3777e+06, 6.3777e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 6.3778e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 6.3779e+06, 
    6.3779e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 6.3782e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 
    6.3784e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3786e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.3789e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3786e+06, 6.3786e+06, 6.3786e+06, 
    6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3785e+06, 6.3784e+06, 
    6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 6.3784e+06, 
    6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3783e+06, 6.3782e+06, 
    6.3782e+06, 6.3782e+06, 6.3782e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3781e+06, 6.3781e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 6.378e+06, 
    6.378e+06, 6.378e+06, 6.378e+06, 6.3781e+06, 6.3781e+06, 6.3781e+06, 
    6.3782e+06, 6.3782e+06, 6.3783e+06, 6.3783e+06, 6.3784e+06, 6.3784e+06, 
    6.3785e+06, 6.3785e+06, 6.3786e+06, 6.3787e+06, 6.3787e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 
    6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 6.3787e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 
    6.3789e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.3788e+06, 
    6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 6.3788e+06, 
    6.3788e+06, 6.3789e+06, 6.3789e+06, 6.3789e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 
    6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.379e+06, 6.379e+06, 6.379e+06, 6.379e+06, 
    6.379e+06, 6.379e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 6.3791e+06, 
    6.3791e+06, 6.3791e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 6.3792e+06, 
    6.3792e+06, 6.3792e+06, 6.3793e+06, 6.3793e+06, 6.3793e+06, 6.3794e+06, 
    6.3794e+06, 6.3794e+06, 6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3796e+06, 
    6.3796e+06, 6.3796e+06, 6.3797e+06, 6.3797e+06, 6.3798e+06, 6.3798e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.38e+06, 
    6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 6.38e+06, 
    6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3799e+06, 6.3798e+06, 6.3798e+06, 
    6.3798e+06, 6.3798e+06, 6.3797e+06, 6.3797e+06, 6.3796e+06, 6.3796e+06, 
    6.3795e+06, 6.3795e+06, 6.3795e+06, 6.3794e+06, 6.3794e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3805e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 
    6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3804e+06, 6.3805e+06, 6.3805e+06, 
    6.3805e+06, 6.3805e+06, 6.3805e+06, 6.3806e+06, 6.3806e+06, 6.3806e+06, 
    6.3807e+06, 6.3807e+06, 6.3807e+06, 6.3808e+06, 6.3808e+06, 6.3808e+06, 
    6.3809e+06, 6.3809e+06, 6.3809e+06, 6.381e+06, 6.381e+06, 6.381e+06, 
    6.381e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3811e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 6.3812e+06, 
    6.3812e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 
    6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3813e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 6.3814e+06, 
    6.3814e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 6.3815e+06, 
    6.3815e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 6.3816e+06, 
    6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 6.3817e+06, 
    6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 6.3818e+06, 
    6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 6.3819e+06, 
    6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 6.382e+06, 
    6.382e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 6.3821e+06, 
    6.3821e+06, 6.3821e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 
    6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3822e+06, 6.3823e+06, 6.3823e+06, 
    6.3823e+06, 6.3823e+06, 6.3823e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 
    6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3824e+06, 6.3825e+06, 6.3825e+06, 
    6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 6.3825e+06, 
    6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3826e+06, 6.3827e+06, 
    6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3827e+06, 6.3828e+06, 6.3828e+06, 
    6.3828e+06, 6.3828e+06, 6.3828e+06, 6.3829e+06, 6.3829e+06, 6.3829e+06, 
    6.3829e+06, 6.3829e+06, 6.383e+06, 6.383e+06, 6.383e+06, 6.383e+06, 
    6.383e+06, 6.383e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 6.3831e+06, 
    6.3831e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3832e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 6.3833e+06, 
    6.3833e+06, 6.3833e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 
    6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3834e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 6.3835e+06, 
    6.3835e+06, 6.3835e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 
    6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3836e+06, 6.3837e+06, 
    6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3837e+06, 6.3838e+06, 
    6.3838e+06, 6.3838e+06, 6.3838e+06, 6.3839e+06, 6.3839e+06, 6.3839e+06, 
    6.3839e+06, 6.3839e+06, 6.3839e+06, 6.384e+06, 6.384e+06, 6.384e+06, 
    6.384e+06, 6.384e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 6.3841e+06, 
    6.3841e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3842e+06, 6.3843e+06, 
    6.3843e+06, 6.3843e+06, 6.3843e+06, 6.3844e+06, 6.3844e+06, 6.3844e+06, 
    6.3844e+06, 6.3845e+06, 6.3845e+06, 6.3845e+06, 6.3846e+06, 6.3846e+06, 
    6.3846e+06, 6.3846e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 6.3847e+06, 
    6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3848e+06, 6.3849e+06, 
    6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.3849e+06, 6.385e+06, 
    6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 6.385e+06, 
    6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 6.3851e+06, 
    6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3852e+06, 6.3853e+06, 
    6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3853e+06, 6.3854e+06, 
    6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3854e+06, 6.3855e+06, 6.3855e+06, 
    6.3855e+06, 6.3855e+06, 6.3855e+06, 6.3856e+06, 6.3856e+06, 6.3856e+06, 
    6.3856e+06, 6.3856e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 6.3857e+06, 
    6.3857e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3858e+06, 6.3859e+06, 
    6.3859e+06, 6.3859e+06, 6.3859e+06, 6.3859e+06, 6.386e+06, 6.386e+06, 
    6.386e+06, 6.386e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 6.3861e+06, 
    6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3862e+06, 6.3863e+06, 6.3863e+06, 
    6.3863e+06, 6.3863e+06, 6.3863e+06, 6.3864e+06, 6.3864e+06, 6.3864e+06, 
    6.3864e+06, 6.3864e+06, 6.3864e+06, 6.3865e+06, 6.3865e+06, 6.3865e+06, 
    6.3865e+06, 6.3865e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 6.3866e+06, 
    6.3867e+06, 6.3867e+06, 6.3867e+06, 6.3868e+06, 6.3868e+06, 6.3868e+06, 
    6.3869e+06, 6.3869e+06, 6.3869e+06, 6.387e+06, 6.387e+06, 6.3871e+06, 
    6.3871e+06, 6.3871e+06, 6.3872e+06, 6.3872e+06, 6.3872e+06, 6.3873e+06, 
    6.3873e+06, 6.3873e+06, 6.3874e+06, 6.3874e+06, 6.3874e+06, 6.3875e+06, 
    6.3875e+06, 6.3875e+06, 6.3875e+06, 6.3876e+06, 6.3876e+06, 6.3876e+06, 
    6.3876e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 6.3877e+06, 
    6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 6.3878e+06, 
    6.3878e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 6.3879e+06, 
    6.3879e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 6.388e+06, 
    6.388e+06, 6.388e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 
    6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3881e+06, 6.3882e+06, 6.3882e+06, 
    6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3882e+06, 6.3883e+06, 
    6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 6.3883e+06, 
    6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 6.3884e+06, 
    6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 6.3885e+06, 
    6.3885e+06, 6.3885e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 
    6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3886e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 6.3887e+06, 
    6.3887e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 6.3888e+06, 
    6.3888e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 6.3889e+06, 
    6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.389e+06, 6.3891e+06, 
    6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3891e+06, 6.3892e+06, 6.3892e+06, 
    6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3892e+06, 6.3893e+06, 
    6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 6.3893e+06, 
    6.3893e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 6.3894e+06, 
    6.3894e+06, 6.3894e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 6.3895e+06, 
    6.3895e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3896e+06, 6.3897e+06, 
    6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3897e+06, 6.3898e+06, 6.3898e+06, 
    6.3898e+06, 6.3898e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 6.3899e+06, 
    6.3899e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.39e+06, 6.3901e+06, 
    6.3901e+06, 6.3901e+06, 6.3901e+06, 6.3902e+06, 6.3902e+06, 6.3902e+06, 
    6.3902e+06, 6.3902e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 6.3903e+06, 
    6.3903e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 6.3904e+06, 
    6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3905e+06, 6.3906e+06, 6.3906e+06, 
    6.3906e+06, 6.3906e+06, 6.3906e+06, 6.3907e+06, 6.3907e+06, 6.3907e+06, 
    6.3907e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 6.3908e+06, 
    6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.3909e+06, 6.391e+06, 
    6.391e+06, 6.391e+06, 6.391e+06, 6.391e+06, 6.3911e+06, 6.3911e+06, 
    6.3911e+06, 6.3911e+06, 6.3911e+06, 6.3912e+06, 6.3912e+06, 6.3912e+06, 
    6.3912e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3913e+06, 6.3914e+06, 
    6.3914e+06, 6.3914e+06, 6.3914e+06, 6.3915e+06, 6.3915e+06, 6.3915e+06, 
    6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3916e+06, 6.3917e+06, 6.3917e+06, 
    6.3917e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3918e+06, 6.3919e+06, 
    6.3919e+06, 6.3919e+06, 6.392e+06, 6.392e+06, 6.392e+06, 6.3921e+06, 
    6.3921e+06, 6.3921e+06, 6.3921e+06, 6.3922e+06, 6.3922e+06, 6.3922e+06, 
    6.3922e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3923e+06, 6.3924e+06, 
    6.3924e+06, 6.3924e+06, 6.3924e+06, 6.3925e+06, 6.3925e+06, 6.3925e+06, 
    6.3925e+06, 6.3926e+06, 6.3926e+06, 6.3926e+06, 6.3927e+06, 6.3927e+06, 
    6.3927e+06, 6.3927e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 6.3928e+06, 
    6.3929e+06, 6.3929e+06, 6.3929e+06, 6.3929e+06, 6.393e+06, 6.393e+06, 
    6.393e+06, 6.393e+06, 6.3931e+06, 6.3931e+06, 6.3931e+06, 6.3932e+06, 
    6.3932e+06, 6.3932e+06, 6.3933e+06, 6.3933e+06, 6.3933e+06, 6.3934e+06, 
    6.3934e+06, 6.3934e+06, 6.3934e+06, 6.3935e+06, 6.3935e+06, 6.3935e+06, 
    6.3936e+06, 6.3936e+06, 6.3936e+06, 6.3937e+06, 6.3937e+06, 6.3937e+06, 
    6.3937e+06, 6.3938e+06, 6.3938e+06, 6.3938e+06, 6.3939e+06, 6.3939e+06, 
    6.3939e+06, 6.3939e+06, 6.394e+06, 6.394e+06, 6.394e+06, 6.394e+06, 
    6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3941e+06, 6.3942e+06, 6.3942e+06, 
    6.3942e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3943e+06, 6.3944e+06, 
    6.3944e+06, 6.3944e+06, 6.3945e+06, 6.3945e+06, 6.3945e+06, 6.3946e+06, 
    6.3946e+06, 6.3946e+06, 6.3947e+06, 6.3947e+06, 6.3948e+06, 6.3948e+06, 
    6.3948e+06, 6.3949e+06, 6.3949e+06, 6.3949e+06, 6.395e+06, 6.395e+06, 
    6.395e+06, 6.3951e+06, 6.3951e+06, 6.3952e+06, 6.3952e+06, 6.3952e+06, 
    6.3953e+06, 6.3953e+06, 6.3953e+06, 6.3954e+06, 6.3954e+06, 6.3955e+06, 
    6.3955e+06, 6.3955e+06, 6.3956e+06, 6.3956e+06, 6.3956e+06, 6.3957e+06, 
    6.3957e+06, 6.3957e+06, 6.3958e+06, 6.3958e+06, 6.3959e+06, 6.3959e+06, 
    6.3959e+06, 6.396e+06, 6.396e+06, 6.396e+06, 6.3961e+06, 6.3961e+06, 
    6.3961e+06, 6.3962e+06, 6.3962e+06, 6.3963e+06, 6.3963e+06, 6.3963e+06, 
    6.3964e+06, 6.3964e+06, 6.3964e+06, 6.3965e+06, 6.3965e+06, 6.3966e+06, 
    6.3966e+06, 6.3966e+06, 6.3967e+06, 6.3967e+06, 6.3967e+06, 6.3968e+06, 
    6.3968e+06, 6.3969e+06, 6.3969e+06, 6.3969e+06, 6.397e+06, 6.397e+06, 
    6.397e+06, 6.3971e+06, 6.3971e+06, 6.3971e+06, 6.3972e+06, 6.3972e+06, 
    6.3973e+06, 6.3973e+06, 6.3973e+06, 6.3974e+06, 6.3974e+06, 6.3974e+06, 
    6.3975e+06, 6.3975e+06, 6.3976e+06, 6.3976e+06, 6.3976e+06, 6.3977e+06, 
    6.3977e+06, 6.3978e+06, 6.3978e+06, 6.3979e+06, 6.3979e+06, 6.3979e+06, 
    6.398e+06, 6.398e+06, 6.3981e+06, 6.3981e+06, 6.3982e+06, 6.3982e+06, 
    6.3983e+06, 6.3983e+06, 6.3984e+06, 6.3984e+06, 6.3985e+06, 6.3985e+06, 
    6.3985e+06, 6.3986e+06, 6.3986e+06, 6.3987e+06, 6.3987e+06, 6.3988e+06, 
    6.3988e+06, 6.3988e+06, 6.3989e+06, 6.3989e+06, 6.399e+06, 6.399e+06, 
    6.399e+06, 6.3991e+06, 6.3991e+06, 6.3992e+06, 6.3992e+06, 6.3992e+06, 
    6.3993e+06, 6.3993e+06, 6.3994e+06, 6.3994e+06, 6.3994e+06, 6.3995e+06, 
    6.3995e+06, 6.3996e+06, 6.3996e+06, 6.3996e+06, 6.3997e+06, 6.3997e+06, 
    6.3997e+06, 6.3998e+06, 6.3998e+06, 6.3999e+06, 6.3999e+06, 6.4e+06, 
    6.4e+06, 6.4e+06, 6.4001e+06, 6.4001e+06, 6.4002e+06, 6.4002e+06, 
    6.4003e+06, 6.4003e+06, 6.4004e+06, 6.4004e+06, 6.4005e+06, 6.4005e+06, 
    6.4006e+06, 6.4006e+06, 6.4007e+06, 6.4007e+06, 6.4008e+06, 6.4008e+06, 
    6.4008e+06, 6.4009e+06, 6.4009e+06, 6.401e+06, 6.401e+06, 6.4011e+06, 
    6.4011e+06, 6.4012e+06, 6.4012e+06, 6.4013e+06, 6.4013e+06, 6.4013e+06, 
    6.4014e+06, 6.4014e+06, 6.4015e+06, 6.4015e+06, 6.4016e+06, 6.4016e+06, 
    6.4017e+06, 6.4017e+06, 6.4018e+06, 6.4018e+06, 6.4019e+06, 6.4019e+06, 
    6.402e+06, 6.402e+06, 6.4021e+06, 6.4021e+06, 6.4021e+06, 6.4022e+06, 
    6.4022e+06, 6.4023e+06, 6.4023e+06, 6.4024e+06, 6.4025e+06, 6.4025e+06, 
    6.4026e+06, 6.4026e+06, 6.4027e+06, 6.4027e+06, 6.4028e+06, 6.4028e+06, 
    6.4029e+06, 6.4029e+06, 6.403e+06, 6.403e+06, 6.403e+06, 6.4031e+06, 
    6.4031e+06, 6.4032e+06, 6.4032e+06, 6.4033e+06, 6.4033e+06, 6.4034e+06, 
    6.4034e+06, 6.4035e+06, 6.4035e+06, 6.4036e+06, 6.4036e+06, 6.4037e+06, 
    6.4037e+06, 6.4038e+06, 6.4038e+06, 6.4039e+06, 6.4039e+06, 6.404e+06, 
    6.404e+06, 6.4041e+06, 6.4041e+06, 6.4042e+06, 6.4042e+06, 6.4043e+06, 
    6.4044e+06, 6.4044e+06, 6.4045e+06, 6.4045e+06, 6.4046e+06, 6.4046e+06, 
    6.4047e+06, 6.4047e+06, 6.4048e+06, 6.4048e+06, 6.4049e+06, 6.4049e+06, 
    6.405e+06, 6.405e+06, 6.4051e+06, 6.4051e+06, 6.4052e+06, 6.4053e+06, 
    6.4053e+06, 6.4054e+06, 6.4054e+06, 6.4055e+06, 6.4055e+06, 6.4056e+06, 
    6.4056e+06, 6.4057e+06, 6.4057e+06, 6.4058e+06, 6.4058e+06, 6.4059e+06, 
    6.406e+06, 6.406e+06, 6.4061e+06, 6.4061e+06, 6.4062e+06, 6.4062e+06, 
    6.4063e+06, 6.4063e+06, 6.4064e+06, 6.4064e+06, 6.4065e+06, 6.4065e+06, 
    6.4066e+06, 6.4066e+06, 6.4067e+06, 6.4067e+06, 6.4068e+06, 6.4068e+06, 
    6.4069e+06, 6.4069e+06, 6.407e+06, 6.407e+06, 6.4071e+06, 6.4071e+06, 
    6.4072e+06, 6.4072e+06, 6.4073e+06, 6.4073e+06, 6.4074e+06, 6.4074e+06, 
    6.4075e+06, 6.4075e+06, 6.4076e+06, 6.4076e+06, 6.4077e+06, 6.4078e+06, 
    6.4078e+06, 6.4079e+06, 6.4079e+06, 6.408e+06, 6.408e+06, 6.4081e+06, 
    6.4082e+06, 6.4082e+06, 6.4083e+06, 6.4083e+06, 6.4084e+06, 6.4084e+06, 
    6.4085e+06, 6.4085e+06, 6.4086e+06, 6.4086e+06, 6.4087e+06, 6.4088e+06, 
    6.4088e+06, 6.4089e+06, 6.4089e+06, 6.409e+06, 6.409e+06, 6.4091e+06, 
    6.4091e+06, 6.4092e+06, 6.4092e+06, 6.4093e+06, 6.4094e+06, 6.4094e+06, 
    6.4095e+06, 6.4095e+06, 6.4096e+06, 6.4096e+06, 6.4097e+06, 6.4097e+06, 
    6.4098e+06, 6.4099e+06, 6.4099e+06, 6.41e+06, 6.41e+06, 6.4101e+06, 
    6.4101e+06, 6.4102e+06, 6.4103e+06, 6.4103e+06, 6.4104e+06, 6.4104e+06, 
    6.4105e+06, 6.4105e+06, 6.4106e+06, 6.4106e+06, 6.4107e+06, 6.4108e+06, 
    6.4108e+06, 6.4109e+06, 6.4109e+06, 6.411e+06, 6.411e+06, 6.4111e+06, 
    6.4111e+06, 6.4112e+06, 6.4112e+06, 6.4113e+06, 6.4114e+06, 6.4114e+06, 
    6.4115e+06, 6.4115e+06, 6.4116e+06, 6.4116e+06, 6.4117e+06, 6.4117e+06, 
    6.4118e+06, 6.4119e+06, 6.4119e+06, 6.412e+06, 6.412e+06, 6.4121e+06, 
    6.4121e+06, 6.4122e+06, 6.4123e+06, 6.4123e+06, 6.4124e+06, 6.4124e+06, 
    6.4125e+06, 6.4125e+06, 6.4126e+06, 6.4126e+06, 6.4127e+06, 6.4128e+06, 
    6.4128e+06, 6.4129e+06, 6.4129e+06, 6.413e+06, 6.413e+06, 6.4131e+06, 
    6.4131e+06, 6.4132e+06, 6.4133e+06, 6.4133e+06, 6.4134e+06, 6.4134e+06, 
    6.4135e+06, 6.4135e+06, 6.4136e+06, 6.4136e+06, 6.4137e+06, 6.4138e+06, 
    6.4138e+06, 6.4139e+06, 6.4139e+06, 6.414e+06, 6.414e+06, 6.4141e+06, 
    6.4141e+06, 6.4142e+06, 6.4143e+06, 6.4143e+06, 6.4144e+06, 6.4144e+06, 
    6.4145e+06, 6.4145e+06, 6.4146e+06, 6.4147e+06, 6.4147e+06, 6.4148e+06, 
    6.4148e+06, 6.4149e+06, 6.415e+06, 6.415e+06, 6.4151e+06, 6.4151e+06, 
    6.4152e+06, 6.4153e+06, 6.4153e+06, 6.4154e+06, 6.4154e+06, 6.4155e+06, 
    6.4156e+06, 6.4156e+06, 6.4157e+06, 6.4157e+06, 6.4158e+06, 6.4159e+06, 
    6.4159e+06, 6.416e+06, 6.416e+06, 6.4161e+06, 6.4161e+06, 6.4162e+06, 
    6.4163e+06, 6.4163e+06, 6.4164e+06, 6.4164e+06, 6.4165e+06, 6.4165e+06, 
    6.4166e+06, 6.4166e+06, 6.4167e+06, 6.4168e+06, 6.4168e+06, 6.4169e+06, 
    6.4169e+06, 6.417e+06, 6.417e+06, 6.4171e+06, 6.4171e+06, 6.4172e+06, 
    6.4172e+06, 6.4173e+06, 6.4174e+06, 6.4174e+06, 6.4175e+06, 6.4175e+06, 
    6.4176e+06, 6.4176e+06, 6.4177e+06, 6.4178e+06, 6.4178e+06, 6.4179e+06, 
    6.4179e+06, 6.418e+06, 6.418e+06, 6.4181e+06, 6.4182e+06, 6.4182e+06, 
    6.4183e+06, 6.4183e+06, 6.4184e+06, 6.4184e+06, 6.4185e+06, 6.4186e+06, 
    6.4186e+06, 6.4187e+06, 6.4187e+06, 6.4188e+06, 6.4188e+06, 6.4189e+06, 
    6.419e+06, 6.419e+06, 6.4191e+06, 6.4191e+06, 6.4192e+06, 6.4192e+06, 
    6.4193e+06, 6.4194e+06, 6.4194e+06, 6.4195e+06, 6.4195e+06, 6.4196e+06, 
    6.4197e+06, 6.4197e+06, 6.4198e+06, 6.4198e+06, 6.4199e+06, 6.42e+06, 
    6.42e+06, 6.4201e+06, 6.4201e+06, 6.4202e+06, 6.4202e+06, 6.4203e+06, 
    6.4204e+06, 6.4204e+06, 6.4205e+06, 6.4205e+06, 6.4206e+06, 6.4207e+06, 
    6.4207e+06, 6.4208e+06, 6.4208e+06, 6.4209e+06, 6.421e+06, 6.421e+06, 
    6.4211e+06, 6.4211e+06, 6.4212e+06, 6.4212e+06, 6.4213e+06, 6.4214e+06, 
    6.4214e+06, 6.4215e+06, 6.4215e+06, 6.4216e+06, 6.4216e+06, 6.4217e+06, 
    6.4218e+06, 6.4218e+06, 6.4219e+06, 6.4219e+06, 6.422e+06, 6.4221e+06, 
    6.4221e+06, 6.4222e+06, 6.4222e+06, 6.4223e+06, 6.4224e+06, 6.4224e+06, 
    6.4225e+06, 6.4226e+06, 6.4226e+06, 6.4227e+06, 6.4227e+06, 6.4228e+06, 
    6.4229e+06, 6.4229e+06, 6.423e+06, 6.4231e+06, 6.4231e+06, 6.4232e+06, 
    6.4232e+06, 6.4233e+06, 6.4233e+06, 6.4234e+06, 6.4235e+06, 6.4235e+06, 
    6.4236e+06, 6.4236e+06, 6.4237e+06, 6.4237e+06, 6.4238e+06, 6.4238e+06, 
    6.4239e+06, 6.4239e+06, 6.424e+06, 6.424e+06, 6.4241e+06, 6.4241e+06, 
    6.4242e+06, 6.4242e+06, 6.4243e+06, 6.4243e+06, 6.4244e+06, 6.4245e+06, 
    6.4245e+06, 6.4246e+06, 6.4246e+06, 6.4247e+06, 6.4247e+06, 6.4248e+06, 
    6.4249e+06, 6.4249e+06, 6.425e+06, 6.425e+06, 6.4251e+06, 6.4252e+06, 
    6.4252e+06, 6.4253e+06, 6.4254e+06, 6.4254e+06, 6.4255e+06, 6.4255e+06, 
    6.4256e+06, 6.4257e+06, 6.4257e+06, 6.4258e+06, 6.4258e+06, 6.4259e+06, 
    6.426e+06, 6.426e+06, 6.4261e+06, 6.4261e+06, 6.4262e+06, 6.4262e+06, 
    6.4263e+06, 6.4264e+06, 6.4264e+06, 6.4265e+06, 6.4265e+06, 6.4266e+06, 
    6.4266e+06, 6.4267e+06, 6.4268e+06, 6.4268e+06, 6.4269e+06, 6.4269e+06, 
    6.427e+06, 6.427e+06, 6.4271e+06, 6.4272e+06, 6.4272e+06, 6.4273e+06, 
    6.4273e+06, 6.4274e+06, 6.4274e+06, 6.4275e+06, 6.4276e+06, 6.4276e+06, 
    6.4277e+06, 6.4277e+06, 6.4278e+06, 6.4278e+06, 6.4279e+06, 6.428e+06, 
    6.428e+06, 6.4281e+06, 6.4281e+06, 6.4282e+06, 6.4283e+06, 6.4283e+06, 
    6.4284e+06, 6.4284e+06, 6.4285e+06, 6.4286e+06, 6.4286e+06, 6.4287e+06, 
    6.4288e+06, 6.4288e+06, 6.4289e+06, 6.4289e+06, 6.429e+06, 6.4291e+06, 
    6.4291e+06, 6.4292e+06, 6.4292e+06, 6.4293e+06, 6.4293e+06, 6.4294e+06, 
    6.4295e+06, 6.4295e+06, 6.4296e+06, 6.4296e+06, 6.4297e+06, 6.4297e+06, 
    6.4298e+06, 6.4298e+06, 6.4299e+06, 6.43e+06, 6.43e+06, 6.4301e+06, 
    6.4301e+06, 6.4302e+06, 6.4303e+06, 6.4303e+06, 6.4304e+06, 6.4304e+06, 
    6.4305e+06, 6.4306e+06, 6.4306e+06, 6.4307e+06, 6.4307e+06, 6.4308e+06, 
    6.4309e+06, 6.4309e+06, 6.431e+06, 6.431e+06, 6.4311e+06, 6.4312e+06, 
    6.4312e+06, 6.4313e+06, 6.4313e+06, 6.4314e+06, 6.4314e+06, 6.4315e+06, 
    6.4316e+06, 6.4316e+06, 6.4317e+06, 6.4317e+06, 6.4318e+06, 6.4318e+06, 
    6.4319e+06, 6.4319e+06, 6.432e+06, 6.432e+06, 6.4321e+06, 6.4322e+06, 
    6.4322e+06, 6.4323e+06, 6.4323e+06, 6.4324e+06, 6.4324e+06, 6.4325e+06, 
    6.4326e+06, 6.4326e+06, 6.4327e+06, 6.4327e+06, 6.4328e+06, 6.4328e+06, 
    6.4329e+06, 6.433e+06, 6.433e+06, 6.4331e+06, 6.4331e+06, 6.4332e+06, 
    6.4333e+06, 6.4333e+06, 6.4334e+06, 6.4334e+06, 6.4335e+06, 6.4336e+06, 
    6.4336e+06, 6.4337e+06, 6.4337e+06, 6.4338e+06, 6.4339e+06, 6.4339e+06, 
    6.434e+06, 6.434e+06, 6.4341e+06, 6.4341e+06, 6.4342e+06, 6.4343e+06, 
    6.4343e+06, 6.4344e+06, 6.4344e+06, 6.4345e+06, 6.4345e+06, 6.4346e+06, 
    6.4347e+06, 6.4347e+06, 6.4348e+06, 6.4348e+06, 6.4349e+06, 6.4349e+06, 
    6.435e+06, 6.4351e+06, 6.4351e+06, 6.4352e+06, 6.4352e+06, 6.4353e+06, 
    6.4354e+06, 6.4354e+06, 6.4355e+06, 6.4355e+06, 6.4356e+06, 6.4357e+06, 
    6.4357e+06, 6.4358e+06, 6.4359e+06, 6.4359e+06, 6.436e+06, 6.436e+06, 
    6.4361e+06, 6.4362e+06, 6.4362e+06, 6.4363e+06, 6.4364e+06, 6.4364e+06, 
    6.4365e+06, 6.4365e+06, 6.4366e+06, 6.4367e+06, 6.4367e+06, 6.4368e+06, 
    6.4368e+06, 6.4369e+06, 6.437e+06, 6.437e+06, 6.4371e+06, 6.4371e+06, 
    6.4372e+06, 6.4372e+06, 6.4373e+06, 6.4373e+06, 6.4374e+06, 6.4374e+06, 
    6.4375e+06, 6.4375e+06, 6.4376e+06, 6.4376e+06, 6.4377e+06, 6.4378e+06, 
    6.4378e+06, 6.4379e+06, 6.4379e+06, 6.438e+06, 6.438e+06, 6.4381e+06, 
    6.4382e+06, 6.4382e+06, 6.4383e+06, 6.4383e+06, 6.4384e+06, 6.4384e+06, 
    6.4385e+06, 6.4386e+06, 6.4386e+06, 6.4387e+06, 6.4387e+06, 6.4388e+06, 
    6.4389e+06, 6.4389e+06, 6.439e+06, 6.439e+06, 6.4391e+06, 6.4392e+06, 
    6.4392e+06, 6.4393e+06, 6.4393e+06, 6.4394e+06, 6.4395e+06, 6.4395e+06, 
    6.4396e+06, 6.4396e+06, 6.4397e+06, 6.4398e+06, 6.4398e+06, 6.4399e+06, 
    6.4399e+06, 6.44e+06, 6.44e+06, 6.4401e+06, 6.4401e+06, 6.4402e+06, 
    6.4402e+06, 6.4403e+06, 6.4403e+06, 6.4404e+06, 6.4405e+06, 6.4405e+06, 
    6.4406e+06, 6.4406e+06, 6.4407e+06, 6.4407e+06, 6.4408e+06, 6.4409e+06, 
    6.4409e+06, 6.441e+06, 6.441e+06, 6.4411e+06, 6.4411e+06, 6.4412e+06, 
    6.4413e+06, 6.4413e+06, 6.4414e+06, 6.4414e+06, 6.4415e+06, 6.4416e+06, 
    6.4416e+06, 6.4417e+06, 6.4418e+06, 6.4418e+06, 6.4419e+06, 6.4419e+06, 
    6.442e+06, 6.4421e+06, 6.4421e+06, 6.4422e+06, 6.4422e+06, 6.4423e+06, 
    6.4423e+06, 6.4424e+06, 6.4425e+06, 6.4425e+06, 6.4426e+06, 6.4426e+06, 
    6.4427e+06, 6.4428e+06, 6.4428e+06, 6.4429e+06, 6.4429e+06, 6.443e+06, 
    6.4431e+06, 6.4431e+06, 6.4432e+06, 6.4432e+06, 6.4433e+06, 6.4434e+06, 
    6.4434e+06, 6.4435e+06, 6.4435e+06, 6.4436e+06, 6.4437e+06, 6.4437e+06, 
    6.4438e+06, 6.4438e+06, 6.4439e+06, 6.4439e+06, 6.444e+06, 6.444e+06, 
    6.4441e+06, 6.4441e+06, 6.4442e+06, 6.4443e+06, 6.4443e+06, 6.4444e+06, 
    6.4444e+06, 6.4445e+06, 6.4445e+06, 6.4446e+06, 6.4446e+06, 6.4447e+06, 
    6.4447e+06, 6.4448e+06, 6.4449e+06, 6.4449e+06, 6.445e+06, 6.445e+06, 
    6.4451e+06, 6.4452e+06, 6.4452e+06, 6.4453e+06, 6.4453e+06, 6.4454e+06, 
    6.4455e+06, 6.4455e+06, 6.4456e+06, 6.4457e+06, 6.4457e+06, 6.4458e+06, 
    6.4458e+06, 6.4459e+06, 6.4459e+06, 6.446e+06, 6.4461e+06, 6.4461e+06, 
    6.4462e+06, 6.4462e+06, 6.4463e+06, 6.4463e+06, 6.4464e+06, 6.4465e+06, 
    6.4465e+06, 6.4466e+06, 6.4466e+06, 6.4467e+06, 6.4467e+06, 6.4468e+06, 
    6.4468e+06, 6.4469e+06, 6.447e+06, 6.447e+06, 6.4471e+06, 6.4471e+06, 
    6.4472e+06, 6.4472e+06, 6.4473e+06, 6.4474e+06, 6.4474e+06, 6.4475e+06, 
    6.4475e+06, 6.4476e+06, 6.4477e+06, 6.4477e+06, 6.4478e+06, 6.4478e+06, 
    6.4479e+06, 6.448e+06, 6.448e+06, 6.4481e+06, 6.4481e+06, 6.4482e+06, 
    6.4482e+06, 6.4483e+06, 6.4484e+06, 6.4484e+06, 6.4485e+06, 6.4485e+06, 
    6.4486e+06, 6.4486e+06, 6.4487e+06, 6.4487e+06, 6.4488e+06, 6.4489e+06, 
    6.4489e+06, 6.449e+06, 6.449e+06, 6.4491e+06, 6.4492e+06, 6.4492e+06, 
    6.4493e+06, 6.4493e+06, 6.4494e+06, 6.4494e+06, 6.4495e+06, 6.4496e+06, 
    6.4496e+06, 6.4497e+06, 6.4497e+06, 6.4498e+06, 6.4499e+06, 6.4499e+06, 
    6.45e+06, 6.45e+06, 6.4501e+06, 6.4502e+06, 6.4502e+06, 6.4503e+06, 
    6.4503e+06, 6.4504e+06, 6.4504e+06, 6.4505e+06, 6.4506e+06, 6.4506e+06, 
    6.4507e+06, 6.4507e+06, 6.4508e+06, 6.4508e+06, 6.4509e+06, 6.451e+06, 
    6.451e+06, 6.4511e+06, 6.4511e+06, 6.4512e+06, 6.4513e+06, 6.4513e+06, 
    6.4514e+06, 6.4514e+06, 6.4515e+06, 6.4516e+06, 6.4516e+06, 6.4517e+06, 
    6.4517e+06, 6.4518e+06, 6.4518e+06, 6.4519e+06, 6.452e+06, 6.452e+06, 
    6.4521e+06, 6.4521e+06, 6.4522e+06, 6.4522e+06, 6.4523e+06, 6.4524e+06, 
    6.4524e+06, 6.4525e+06, 6.4525e+06, 6.4526e+06, 6.4526e+06, 6.4527e+06, 
    6.4527e+06, 6.4528e+06, 6.4529e+06, 6.4529e+06, 6.453e+06, 6.453e+06, 
    6.4531e+06, 6.4532e+06, 6.4532e+06, 6.4533e+06, 6.4533e+06, 6.4534e+06, 
    6.4535e+06, 6.4535e+06, 6.4536e+06, 6.4536e+06, 6.4537e+06, 6.4538e+06, 
    6.4538e+06, 6.4539e+06, 6.4539e+06, 6.454e+06, 6.454e+06, 6.4541e+06, 
    6.4541e+06, 6.4542e+06, 6.4543e+06, 6.4543e+06, 6.4544e+06, 6.4544e+06, 
    6.4545e+06, 6.4545e+06, 6.4546e+06, 6.4546e+06, 6.4547e+06, 6.4547e+06, 
    6.4548e+06, 6.4548e+06, 6.4549e+06, 6.455e+06, 6.455e+06, 6.4551e+06, 
    6.4551e+06, 6.4552e+06, 6.4552e+06, 6.4553e+06, 6.4554e+06, 6.4554e+06, 
    6.4555e+06, 6.4555e+06, 6.4556e+06, 6.4557e+06, 6.4557e+06, 6.4558e+06, 
    6.4559e+06, 6.4559e+06, 6.456e+06, 6.456e+06, 6.4561e+06, 6.4562e+06, 
    6.4562e+06, 6.4563e+06, 6.4563e+06, 6.4564e+06, 6.4565e+06, 6.4565e+06, 
    6.4566e+06, 6.4566e+06, 6.4567e+06, 6.4567e+06, 6.4568e+06, 6.4568e+06, 
    6.4569e+06 ;

 impact_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1 =
  0.022189, 0.02217, 0.022151, 0.02213, 0.022112, 0.022093, 0.022075, 
    0.022057, 0.022038, 0.022019, 0.022001, 0.021982, 0.021963, 0.021943, 
    0.021921, 0.021901, 0.02188, 0.021858, 0.021834, 0.021811, 0.021787, 
    0.021764, 0.021742, 0.021721, 0.021699, 0.021677, 0.021656, 0.021633, 
    0.021609, 0.021586, 0.021564, 0.021544, 0.021525, 0.021508, 0.021492, 
    0.021478, 0.021466, 0.021454, 0.021441, 0.021427, 0.021415, 0.021403, 
    0.021393, 0.021383, 0.021375, 0.021369, 0.021364, 0.021358, 0.021352, 
    0.021346, 0.02134, 0.021334, 0.021329, 0.021324, 0.021318, 0.021312, 
    0.021305, 0.021297, 0.021288, 0.021278, 0.021269, 0.021259, 0.021249, 
    0.021237, 0.021224, 0.02121, 0.021195, 0.021178, 0.021158, 0.021142, 
    0.021124, 0.021105, 0.021087, 0.021069, 0.021051, 0.021033, 0.021017, 
    0.021, 0.020983, 0.020965, 0.020948, 0.020931, 0.020913, 0.020897, 
    0.020882, 0.020863, 0.020845, 0.020827, 0.020808, 0.020791, 0.020769, 
    0.020749, 0.020729, 0.020709, 0.020688, 0.020674, 0.020659, 0.020647, 
    0.020636, 0.020621, 0.02061, 0.020598, 0.020587, 0.020577, 0.020568, 
    0.020557, 0.020553, 0.020547, 0.020541, 0.020535, 0.020524, 0.020517, 
    0.02051, 0.020504, 0.020498, 0.020491, 0.020484, 0.020476, 0.020468, 
    0.020461, 0.020449, 0.020437, 0.020425, 0.020413, 0.020399, 0.020385, 
    0.02037, 0.020355, 0.020339, 0.020319, 0.020301, 0.020282, 0.02026, 
    0.020235, 0.020209, 0.020181, 0.020153, 0.020123, 0.020093, 0.020062, 
    0.020031, 0.019998, 0.019967, 0.019936, 0.019908, 0.01988, 0.019851, 
    0.019822, 0.019791, 0.01976, 0.019734, 0.019706, 0.019679, 0.019652, 
    0.019623, 0.019593, 0.019568, 0.019544, 0.01952, 0.019498, 0.019471, 
    0.019447, 0.019421, 0.019395, 0.019369, 0.019342, 0.019312, 0.019285, 
    0.019257, 0.019229, 0.019201, 0.01917, 0.019143, 0.019117, 0.019091, 
    0.019065, 0.01904, 0.019015, 0.018991, 0.018966, 0.018947, 0.018925, 
    0.018903, 0.018883, 0.018863, 0.018844, 0.018828, 0.018809, 0.018794, 
    0.018783, 0.018775, 0.018768, 0.018762, 0.018755, 0.018752, 0.018751, 
    0.018748, 0.018746, 0.018745, 0.018746, 0.018746, 0.018748, 0.018744, 
    0.018742, 0.01874, 0.018736, 0.018732, 0.018728, 0.018725, 0.01872, 
    0.018711, 0.018701, 0.018692, 0.018683, 0.018672, 0.018658, 0.018645, 
    0.018626, 0.018609, 0.018591, 0.018575, 0.018559, 0.018541, 0.018522, 
    0.018501, 0.018479, 0.018454, 0.018434, 0.018412, 0.018385, 0.018357, 
    0.018327, 0.018296, 0.018265, 0.018238, 0.01821, 0.01818, 0.01815, 
    0.018119, 0.018087, 0.018055, 0.018027, 0.018001, 0.017975, 0.017949, 
    0.017923, 0.017897, 0.017873, 0.017845, 0.017815, 0.017787, 0.017761, 
    0.017735, 0.017712, 0.017685, 0.017663, 0.017641, 0.017617, 0.017595, 
    0.017576, 0.017561, 0.017546, 0.017534, 0.017518, 0.017505, 0.017493, 
    0.017478, 0.01746, 0.017441, 0.017422, 0.017402, 0.017379, 0.017357, 
    0.017335, 0.017314, 0.017294, 0.017274, 0.017256, 0.017233, 0.017211, 
    0.01719, 0.017171, 0.017156, 0.017142, 0.017129, 0.017116, 0.017103, 
    0.017088, 0.017078, 0.01707, 0.017058, 0.017046, 0.017035, 0.017025, 
    0.017012, 0.017006, 0.016999, 0.016991, 0.016981, 0.016967, 0.016949, 
    0.016928, 0.016907, 0.016884, 0.016861, 0.016836, 0.01681, 0.016784, 
    0.016761, 0.016737, 0.016709, 0.016683, 0.01666, 0.016635, 0.01661, 
    0.016583, 0.016557, 0.016528, 0.016497, 0.016465, 0.016434, 0.016404, 
    0.016375, 0.016346, 0.016318, 0.016291, 0.016269, 0.016249, 0.016231, 
    0.016215, 0.016201, 0.016189, 0.016178, 0.016169, 0.016161, 0.016153, 
    0.016146, 0.016139, 0.016132, 0.016123, 0.016114, 0.016104, 0.016092, 
    0.016081, 0.016071, 0.016061, 0.016048, 0.016032, 0.016015, 0.015996, 
    0.015977, 0.01596, 0.01594, 0.015918, 0.015895, 0.015871, 0.015848, 
    0.015826, 0.015803, 0.01578, 0.015756, 0.015731, 0.015707, 0.015683, 
    0.015659, 0.015634, 0.015607, 0.015578, 0.015546, 0.01552, 0.015493, 
    0.015461, 0.01543, 0.015405, 0.015382, 0.01536, 0.015338, 0.015318, 
    0.015301, 0.015283, 0.015265, 0.015249, 0.015232, 0.015217, 0.015201, 
    0.015188, 0.015176, 0.015164, 0.015151, 0.015135, 0.015121, 0.015108, 
    0.015096, 0.015081, 0.015072, 0.015063, 0.015056, 0.015046, 0.015037, 
    0.015029, 0.015022, 0.015013, 0.015007, 0.015002, 0.014998, 0.014991, 
    0.014987, 0.014982, 0.014974, 0.014964, 0.014948, 0.014932, 0.014918, 
    0.014903, 0.014886, 0.014868, 0.01485, 0.014831, 0.014812, 0.014789, 
    0.014765, 0.014739, 0.014712, 0.014682, 0.014653, 0.014623, 0.014596, 
    0.014565, 0.014532, 0.014495, 0.014464, 0.01443, 0.014396, 0.014359, 
    0.014325, 0.014293, 0.014263, 0.014235, 0.011673, 0.011652, 0.011632, 
    0.011613, 0.011593, 0.011575, 0.011552, 0.011538, 0.011516, 0.011496, 
    0.011476, 0.011457, 0.011434, 0.011414, 0.011395, 0.011374, 0.01135, 
    0.011328, 0.01131, 0.011284, 0.011259, 0.011234, 0.01121, 0.011188, 
    0.011165, 0.011144, 0.011123, 0.011103, 0.011085, 0.011066, 0.011048, 
    0.011031, 0.011018, 0.011003, 0.010989, 0.010973, 0.01096, 0.010948, 
    0.010936, 0.010923, 0.010912, 0.010902, 0.010893, 0.010884, 0.010876, 
    0.010864, 0.010856, 0.010848, 0.01084, 0.010832, 0.010826, 0.010818, 
    0.010805, 0.010791, 0.010779, 0.010768, 0.010757, 0.010745, 0.010733, 
    0.010719, 0.010705, 0.010689, 0.010673, 0.010656, 0.010638, 0.010621, 
    0.010604, 0.010582, 0.010566, 0.010547, 0.010528, 0.01051, 0.010492, 
    0.010474, 0.010456, 0.010439, 0.010422, 0.010405, 0.010388, 0.010377, 
    0.01036, 0.010343, 0.010325, 0.010308, 0.010291, 0.010274, 0.010258, 
    0.010242, 0.010226, 0.01021, 0.010194, 0.010178, 0.010162, 0.010147, 
    0.010133, 0.010119, 0.010106, 0.010092, 0.010078, 0.010064, 0.010049, 
    0.010035, 0.010021, 0.010007, 0.0099935, 0.0099806, 0.0099633, 0.0099479, 
    0.0099327, 0.0099184, 0.0099037, 0.0098904, 0.0098761, 0.0098624, 
    0.0098479, 0.0098332, 0.0098184, 0.009804, 0.0097898, 0.009776, 
    0.0097618, 0.0097473, 0.0097326, 0.0097172, 0.0097021, 0.0096864, 
    0.0096709, 0.0096551, 0.009639, 0.009623, 0.009607, 0.0095912, 0.0095755, 
    0.00956, 0.0095445, 0.0095288, 0.0095129, 0.0094969, 0.0094807, 
    0.0094649, 0.0094491, 0.0094339, 0.0094188, 0.0094044, 0.0093905, 
    0.0093767, 0.0093633, 0.0093495, 0.0093354, 0.0093207, 0.0093058, 
    0.0092902, 0.0092742, 0.0092582, 0.0092421, 0.0092265, 0.0092109, 
    0.0091953, 0.0091797, 0.0091641, 0.0091487, 0.0091333, 0.0091182, 
    0.0091034, 0.009089, 0.0090747, 0.0090606, 0.0090464, 0.0090328, 
    0.0090191, 0.0090064, 0.0089935, 0.0089813, 0.0089684, 0.0089561, 
    0.0089433, 0.0089302, 0.0089169, 0.0089036, 0.0088903, 0.0088771, 
    0.0088627, 0.0088483, 0.0088334, 0.0088182, 0.0088037, 0.0087887, 
    0.0087748, 0.0087607, 0.0087472, 0.008734, 0.0087206, 0.0087075, 
    0.0086945, 0.0086818, 0.0086689, 0.0086559, 0.0086424, 0.0086286, 
    0.008614, 0.0085988, 0.008583, 0.0085664, 0.0085496, 0.0085327, 
    0.0085164, 0.0085003, 0.0084845, 0.0084687, 0.0084527, 0.0084367, 
    0.0084206, 0.0084044, 0.0083881, 0.0083717, 0.0083551, 0.0083384, 
    0.0083216, 0.0083048, 0.0082878, 0.0082711, 0.0082541, 0.008237, 0.00822, 
    0.0082032, 0.0081863, 0.0081695, 0.0081527, 0.0081357, 0.008119, 
    0.0081023, 0.0080857, 0.0080698, 0.0080541, 0.0080389, 0.0080241, 
    0.0080099, 0.0079959, 0.0079823, 0.0079691, 0.0079565, 0.0079446, 
    0.0079316, 0.0079189, 0.0079054, 0.0078913, 0.0078772, 0.0078623, 
    0.0078477, 0.007833, 0.0078182, 0.0078038, 0.0077896, 0.0077755, 
    0.0077617, 0.0077479, 0.0077344, 0.0077212, 0.0077082, 0.0076955, 
    0.007683, 0.0076707, 0.0076585, 0.0076465, 0.0076348, 0.0076233, 
    0.007612, 0.0076008, 0.00759, 0.0075791, 0.0075683, 0.0075574, 0.0075465, 
    0.0075358, 0.0075249, 0.0075141, 0.0075031, 0.0074922, 0.0074809, 
    0.0074694, 0.0074578, 0.0074458, 0.0074333, 0.0074206, 0.0074078, 
    0.0073949, 0.0073817, 0.0073683, 0.0073546, 0.0073404, 0.0073261, 
    0.0073113, 0.0072962, 0.0072811, 0.0072657, 0.0072504, 0.0072353, 
    0.0072201, 0.0072049, 0.0071899, 0.0071749, 0.0071601, 0.0071453, 
    0.0071306, 0.0071162, 0.0071019, 0.0070876, 0.0070734, 0.0070593, 
    0.0070453, 0.0070314, 0.0070176, 0.0070038, 0.0069901, 0.0069766, 
    0.0069629, 0.0069491, 0.0069355, 0.0069219, 0.0069084, 0.0068948, 
    0.0068813, 0.0068677, 0.006854, 0.0068404, 0.0068267, 0.0068131, 
    0.0067995, 0.0067859, 0.0067726, 0.006759, 0.0067455, 0.006732, 
    0.0067185, 0.0067051, 0.0066917, 0.0066784, 0.0066652, 0.0066522, 
    0.0066394, 0.0066266, 0.0066141, 0.0066015, 0.006589, 0.0065768, 
    0.0065646, 0.0065526, 0.0065406, 0.0065287, 0.006517, 0.0065052, 
    0.0064935, 0.0064818, 0.0064699, 0.0064577, 0.0064452, 0.0064326, 
    0.0064198, 0.0064068, 0.0063933, 0.0063798, 0.0063663, 0.0063527, 
    0.0063391, 0.0063254, 0.0063118, 0.0062983, 0.0062847, 0.0062709, 
    0.0062571, 0.0062433, 0.0062297, 0.0062161, 0.0062028, 0.00619, 
    0.0061776, 0.0061659, 0.0061547, 0.0061439, 0.0061336, 0.0061237, 
    0.0061141, 0.0061049, 0.006096, 0.0060872, 0.0060788, 0.0060704, 
    0.0060624, 0.0060544, 0.0060467, 0.0060392, 0.0060315, 0.0060238, 
    0.0060158, 0.0060078, 0.0059994, 0.0059909, 0.0059821, 0.005973, 
    0.0059639, 0.0059546, 0.0059448, 0.0059347, 0.0059242, 0.0059132, 
    0.0059018, 0.00589, 0.0058778, 0.0058654, 0.0058526, 0.0058395, 
    0.0058261, 0.0058125, 0.0057986, 0.0057844, 0.0057699, 0.0057552, 
    0.0057405, 0.0057255, 0.0057103, 0.005695, 0.0056797, 0.0056645, 
    0.0056494, 0.0056343, 0.0056194, 0.0056046, 0.00559, 0.0055753, 
    0.0055606, 0.0055458, 0.0055309, 0.0055158, 0.0055004, 0.0054846, 
    0.0054687, 0.0054528, 0.0054368, 0.0054208, 0.0054048, 0.0053888, 
    0.0053728, 0.0053569, 0.005341, 0.0053254, 0.0053099, 0.0052944, 
    0.005279, 0.0052636, 0.0052484, 0.0052333, 0.0052183, 0.0052034, 
    0.0051886, 0.0051738, 0.005159, 0.0051442, 0.0051293, 0.0051143, 
    0.0050992, 0.0050839, 0.0050687, 0.0050534, 0.005038, 0.0050226, 
    0.0050071, 0.0049914, 0.0049758, 0.0049602, 0.0049447, 0.0049292, 
    0.0049136, 0.0048978, 0.0048817, 0.0048655, 0.004849, 0.0048323, 
    0.0048155, 0.0047987, 0.0047818, 0.0047649, 0.004748, 0.0047314, 
    0.0047149, 0.0046986, 0.0046825, 0.0046666, 0.0046506, 0.0046351, 
    0.0046202, 0.0046054, 0.0045912, 0.0045772, 0.0045633, 0.0045497, 
    0.0045362, 0.004523, 0.00451, 0.0044972, 0.0044843, 0.0044714, 0.0044583, 
    0.004445, 0.0044315, 0.0044176, 0.0044038, 0.0043898, 0.0043756, 
    0.0043612, 0.0043465, 0.0043315, 0.0043165, 0.0043013, 0.0042859, 
    0.0042704, 0.0042549, 0.0042392, 0.0042236, 0.0042081, 0.0041926, 
    0.0041769, 0.0041611, 0.0041453, 0.0041292, 0.0041132, 0.0040972, 
    0.0040813, 0.0040654, 0.0040499, 0.0040347, 0.00402, 0.0040059, 
    0.0039921, 0.0039787, 0.0039655, 0.0039527, 0.0039399, 0.0039273, 
    0.0039148, 0.0039021, 0.0038894, 0.0038768, 0.0038642, 0.0038517, 
    0.0038392, 0.0038268, 0.0038144, 0.0038019, 0.0037891, 0.0037761, 
    0.0037632, 0.0037501, 0.0037372, 0.0037241, 0.0037109, 0.0036977, 
    0.0036845, 0.0036713, 0.0036582, 0.0036453, 0.0036323, 0.0036192, 
    0.0036062, 0.003593, 0.0035799, 0.0035666, 0.0035534, 0.0035403, 
    0.0035273, 0.0035143, 0.0035012, 0.0034881, 0.0034751, 0.0034621, 
    0.0034492, 0.0034364, 0.0034235, 0.0034108, 0.0033982, 0.0033857, 
    0.0033734, 0.0033611, 0.0033487, 0.0033361, 0.0033233, 0.0033105, 
    0.0032976, 0.0032846, 0.0032714, 0.0032579, 0.0032445, 0.003231, 
    0.0032177, 0.0032044, 0.0031911, 0.0031779, 0.0031648, 0.0031516, 
    0.0031386, 0.0031255, 0.0031125, 0.0030995, 0.0030865, 0.0030736, 
    0.0030605, 0.0030475, 0.0030344, 0.0030213, 0.0030082, 0.0029952, 
    0.0029823, 0.0029695, 0.0029568, 0.0029441, 0.0029318, 0.0029195, 
    0.0029074, 0.0028957, 0.0028842, 0.0028731, 0.0028621, 0.0028513, 
    0.0028406, 0.00283, 0.0028194, 0.0028089, 0.0027984, 0.002788, 0.0027777, 
    0.0027673, 0.002757, 0.0027466, 0.0027362, 0.0027258, 0.0027154, 
    0.0027049, 0.0026945, 0.002684, 0.0026736, 0.0026631, 0.0026527, 
    0.0026423, 0.0026319, 0.0026214, 0.0026108, 0.0025999, 0.002589, 
    0.002578, 0.0025669, 0.0025557, 0.0025443, 0.0025328, 0.0025213, 
    0.0025098, 0.0024982, 0.0024867, 0.0024753, 0.0024638, 0.0024523, 
    0.0024408, 0.0024294, 0.0024178, 0.0024063, 0.0023948, 0.0023834, 
    0.002372, 0.0023606, 0.0023493, 0.002338, 0.0023267, 0.0023153, 0.002304, 
    0.0022926, 0.0022812, 0.0022698, 0.0022585, 0.0022472, 0.002236, 
    0.0022249, 0.002214, 0.0022035, 0.0021931, 0.0021828, 0.0021727, 
    0.0021628, 0.002153, 0.0021432, 0.0021335, 0.0021238, 0.0021143, 
    0.0021047, 0.0020951, 0.0020855, 0.0020759, 0.0020662, 0.0020563, 
    0.0020465, 0.0020366, 0.0020267, 0.0020167, 0.0020066, 0.0019967, 
    0.0019867, 0.0019766, 0.0019663, 0.0019559, 0.0019452, 0.0019345, 
    0.0019234, 0.0019124, 0.0019013, 0.0018901, 0.0018789, 0.0018675, 
    0.0018561, 0.0018445, 0.001833, 0.0018215, 0.0018101, 0.0017987, 
    0.0017876, 0.0017766, 0.0017658, 0.0017552, 0.0017448, 0.0017345, 
    0.0017245, 0.0017146, 0.0017049, 0.0016956, 0.0016864, 0.0016775, 
    0.001669, 0.0016606, 0.0016524, 0.0016445, 0.0016366, 0.0016289, 
    0.0016211, 0.0016133, 0.0016056, 0.0015979, 0.0015902, 0.0015825, 
    0.0015749, 0.0015672, 0.0015597, 0.001552, 0.0015444, 0.0015367, 
    0.0015289, 0.0015211, 0.0015134, 0.0015057, 0.0014979, 0.0014901, 
    0.0014822, 0.0014743, 0.0014664, 0.0014584, 0.0014505, 0.0014425, 
    0.0014347, 0.0014268, 0.0014189, 0.0014111, 0.0014033, 0.0013955, 
    0.0013878, 0.0013802, 0.0013725, 0.001365, 0.0013575, 0.0013501, 
    0.0013426, 0.0013352, 0.0013277, 0.0013203, 0.0013128, 0.0013054, 
    0.0012979, 0.0012904, 0.001283, 0.0012756, 0.0012682, 0.0012607, 
    0.0012532, 0.0012456, 0.0012379, 0.0012301, 0.0012223, 0.0012145, 
    0.0012066, 0.0011988, 0.0011909, 0.001183, 0.0011753, 0.0011675, 
    0.0011597, 0.0011519, 0.0011441, 0.0011363, 0.0011285, 0.0011208, 
    0.0011131, 0.0011055, 0.0010979, 0.0010905, 0.0010832, 0.001076, 
    0.001069, 0.001062, 0.0010553, 0.0010486, 0.0010422, 0.0010358, 
    0.0010296, 0.0010235, 0.0010176, 0.0010118, 0.0010063, 0.001001, 
    0.00099604, 0.00099119, 0.00098647, 0.00098178, 0.00097728, 0.00097282, 
    0.00096826, 0.00096376, 0.00095923, 0.00095477, 0.00095022, 0.00094567, 
    0.00094099, 0.00093625, 0.00093145, 0.00092651, 0.00092144, 0.00091617, 
    0.00091076, 0.00090509, 0.00089923, 0.00089331, 0.0008872, 0.0008809, 
    0.00087444, 0.0008678, 0.00086104, 0.0008541, 0.00084703, 0.0008399, 
    0.0008328, 0.00082571, 0.00081859, 0.00081144, 0.00080423, 0.0007971, 
    0.00079003, 0.00078302, 0.00077601, 0.00076906, 0.0007622, 0.00075544, 
    0.00074887, 0.00074239, 0.00073607, 0.0007299, 0.00072392, 0.00071805, 
    0.00071238, 0.00070698, 0.00070178, 0.0006968, 0.0006919, 0.00068724, 
    0.00068277, 0.00067844, 0.00067413, 0.00066991, 0.00066577, 0.00066172, 
    0.00065775, 0.00065381, 0.00064989, 0.00064593, 0.00064191, 0.00063791, 
    0.00063381, 0.00062965, 0.00062542, 0.00062096, 0.00061649, 0.00061182, 
    0.0006071, 0.00060228, 0.00059738, 0.00059249, 0.00058758, 0.00058278, 
    0.00057806, 0.00057342, 0.00056888, 0.00056434, 0.00055988, 0.00055545, 
    0.00055106, 0.00054671, 0.00054239, 0.00053816, 0.00053403, 0.00052994, 
    0.00052584, 0.00052189, 0.00051813, 0.00051448, 0.00051097, 0.00050752, 
    0.00050419, 0.00050102, 0.00049789, 0.00049481, 0.0004918, 0.00048885, 
    0.00048593, 0.00048299, 0.00047999, 0.00047699, 0.00047396, 0.00047093, 
    0.00046784, 0.00046462, 0.00046138, 0.00045808, 0.00045473, 0.00045119, 
    0.0004476, 0.00044395, 0.00044029, 0.0004366, 0.00043286, 0.00042914, 
    0.00042552, 0.00042188, 0.00041838, 0.0004149, 0.00041148, 0.00040824, 
    0.00040504, 0.00040192, 0.00039891, 0.00039599, 0.00039312, 0.00039031, 
    0.00038753, 0.00038479, 0.00038214, 0.0003796, 0.00037703, 0.00037454, 
    0.00037211, 0.00036973, 0.00036749, 0.00036533, 0.0003632, 0.00036104, 
    0.00035887, 0.00035676, 0.0003547, 0.00035265, 0.00035063, 0.00034876, 
    0.00034692, 0.00034506, 0.0003432, 0.00034137, 0.00033951, 0.00033764, 
    0.00033576, 0.00033395, 0.00033212, 0.00033032, 0.00032851, 0.00032677, 
    0.00032504, 0.00032337, 0.00032166, 0.00031986, 0.00031799, 0.00031601, 
    0.00031401, 0.00031188, 0.00030965, 0.00030731, 0.00030488, 0.00030236, 
    0.00029973, 0.00029698, 0.00029414, 0.00029126, 0.00028831, 0.00028526, 
    0.00028213, 0.00027894, 0.00027567, 0.00027248, 0.00026923, 0.00026598, 
    0.00026285, 0.00025971, 0.00025668, 0.00025368, 0.00025074, 0.00024797, 
    0.00024521, 0.00024256, 0.00023997, 0.00023741, 0.00023507, 0.00023281, 
    0.00023072, 0.0002288, 0.00022699, 0.00022539, 0.00022399, 0.00022266, 
    0.00022132, 0.0002201, 0.00021888, 0.00021772, 0.0002166, 0.00021557, 
    0.00021463, 0.00021376, 0.00021289, 0.00021201, 0.00021109, 0.00021009, 
    0.00020896, 0.00020775, 0.00020647, 0.00020509, 0.00020364, 0.00020214, 
    0.00020061, 0.00019905, 0.00019745, 0.00019584, 0.00019419, 0.00019256, 
    0.00019091, 0.0001893, 0.00018772, 0.00018616, 0.00018461, 0.00018313, 
    0.00018166, 0.00018032, 0.00017909, 0.00017793, 0.00017687, 0.00017584, 
    0.00017488, 0.0001739, 0.00017298, 0.00017212, 0.00017132, 0.00017052, 
    0.00016976, 0.00016896, 0.00016816, 0.0001674, 0.00016661, 0.00016573, 
    0.00016488, 0.0001639, 0.00016291, 0.00016179, 0.00016058, 0.00015936, 
    0.00015803, 0.00015671, 0.00015527, 0.00015378, 0.00015224, 0.00015078, 
    0.00014929, 0.00014773, 0.00014618, 0.00014465, 0.00014308, 0.00014155, 
    0.00014007, 0.00013865, 0.00013731, 0.00013601, 0.00013476, 0.00013356, 
    0.00013239, 0.00013132, 0.00013026, 0.00012929, 0.0001284, 0.0001275, 
    0.00012666, 0.00012591, 0.00012517, 0.00012446, 0.00012375, 0.0001231, 
    0.00012244, 0.00012179, 0.0001211, 0.00012042, 0.00011976, 0.000119, 
    0.00011817, 0.00011725, 0.00011618, 0.00011516, 0.00011404, 0.00011286, 
    0.00011168, 0.00011043, 0.00010912, 0.00010779, 0.0001065, 0.0001052, 
    0.0001039, 0.00010261, 0.00010135, 0.00010011, 9.898e-05, 9.7905e-05, 
    9.6851e-05, 9.5872e-05, 9.4819e-05, 9.3797e-05, 9.2714e-05, 9.1686e-05, 
    9.0734e-05, 8.9782e-05, 8.8917e-05, 8.8053e-05, 8.7292e-05, 8.6581e-05, 
    8.5998e-05, 8.5514e-05, 8.5088e-05, 8.4735e-05, 8.4488e-05, 8.431e-05, 
    8.4283e-05, 8.4276e-05, 8.4461e-05, 8.4737e-05, 8.5147e-05, 8.5627e-05, 
    8.6138e-05, 8.6623e-05, 8.7141e-05, 8.7604e-05, 8.8035e-05, 8.8444e-05, 
    8.8792e-05, 8.9085e-05, 8.9297e-05, 8.9339e-05, 8.9287e-05, 8.9025e-05, 
    8.8758e-05, 8.8383e-05, 8.793e-05, 8.742e-05, 8.6878e-05, 8.6327e-05, 
    8.5737e-05, 8.5147e-05, 8.449e-05, 8.3635e-05, 8.2747e-05, 8.1737e-05, 
    8.0595e-05, 7.9486e-05, 7.8216e-05, 7.6924e-05, 7.5585e-05, 7.4195e-05, 
    7.2882e-05, 7.1453e-05, 7.0007e-05, 6.8624e-05, 6.7241e-05, 6.589e-05, 
    6.4563e-05, 6.3325e-05, 6.2242e-05, 6.1237e-05, 6.0312e-05, 5.9501e-05, 
    5.8714e-05, 5.8023e-05, 5.7403e-05, 5.6811e-05, 5.6186e-05, 5.5597e-05, 
    5.5033e-05, 5.4507e-05, 5.4024e-05, 5.3556e-05, 5.3128e-05, 5.2688e-05, 
    5.2159e-05, 5.1628e-05, 5.1018e-05, 5.0352e-05, 4.9658e-05, 4.9021e-05, 
    4.8402e-05, 4.7876e-05, 4.7351e-05, 4.6856e-05, 4.6384e-05, 4.5952e-05, 
    4.5569e-05, 4.5196e-05, 4.4984e-05, 4.4823e-05, 4.471e-05, 4.4688e-05, 
    4.4645e-05, 4.4635e-05, 4.4635e-05, 4.471e-05, 4.4687e-05, 4.4703e-05, 
    4.4719e-05, 4.4769e-05, 4.4875e-05, 4.4914e-05, 4.4909e-05, 4.4977e-05, 
    4.5037e-05, 4.5053e-05, 4.5148e-05, 4.5174e-05, 4.5199e-05, 4.5288e-05, 
    4.5341e-05, 4.5474e-05, 4.5599e-05, 4.5745e-05, 4.5929e-05, 4.6125e-05, 
    4.6259e-05, 4.6239e-05, 4.615e-05, 4.6047e-05, 4.5999e-05, 4.5968e-05, 
    4.6001e-05, 4.5987e-05, 4.5788e-05, 4.5557e-05, 4.5246e-05, 4.4779e-05, 
    4.4261e-05, 4.3713e-05, 4.3152e-05, 4.2571e-05, 4.2138e-05, 4.1787e-05, 
    4.1546e-05, 4.1401e-05, 4.1361e-05, 4.1433e-05, 4.1621e-05, 4.2035e-05, 
    4.2627e-05, 4.3446e-05, 4.449e-05, 4.575e-05, 4.7139e-05, 4.863e-05, 
    5.0205e-05, 5.1828e-05, 5.3408e-05, 5.4959e-05, 5.6418e-05, 5.7816e-05, 
    5.9098e-05, 6.0245e-05, 6.1169e-05, 6.1863e-05, 6.2457e-05, 6.2785e-05, 
    6.2959e-05, 6.3e-05, 6.2789e-05, 6.2447e-05, 6.1804e-05, 6.0923e-05, 
    5.9836e-05, 5.8535e-05, 5.7021e-05, 5.5294e-05, 5.3332e-05, 5.12e-05, 
    4.9038e-05, 4.6736e-05, 4.4393e-05, 4.1994e-05, 3.9615e-05, 3.7196e-05, 
    3.4868e-05, 3.264e-05, 3.0375e-05, 2.8303e-05, 2.6416e-05, 2.4736e-05, 
    2.3378e-05, 2.2441e-05, 2.1756e-05, 2.1212e-05, 2.0982e-05, 2.0907e-05, 
    2.0943e-05, 2.1208e-05, 2.1578e-05, 2.2065e-05, 2.2664e-05, 2.3445e-05, 
    2.4379e-05, 2.5398e-05, 2.6485e-05, 2.7499e-05, 2.8489e-05, 2.9313e-05, 
    3.0188e-05, 3.0942e-05, 3.1696e-05, 3.2403e-05, 3.3072e-05, 3.366e-05, 
    3.4128e-05, 3.4551e-05, 3.4898e-05, 3.5121e-05, 3.5216e-05, 3.5245e-05, 
    3.5159e-05, 3.4919e-05, 3.4536e-05, 3.3996e-05, 3.3327e-05, 3.255e-05, 
    3.1723e-05, 3.0776e-05, 2.9928e-05, 2.8919e-05, 2.8077e-05, 2.7274e-05, 
    2.6531e-05, 2.5889e-05, 2.5287e-05, 2.4773e-05, 2.4293e-05, 2.3868e-05, 
    2.3358e-05, 2.2963e-05, 2.2622e-05, 2.2363e-05, 2.2192e-05, 2.2102e-05, 
    2.1977e-05, 2.191e-05, 2.1872e-05, 2.1736e-05, 2.17e-05, 2.1769e-05, 
    2.1931e-05, 2.2176e-05, 2.2615e-05, 2.3168e-05, 2.3806e-05, 2.4608e-05, 
    2.5596e-05, 2.6692e-05, 2.789e-05, 2.9077e-05, 3.0257e-05, 3.137e-05, 
    3.2505e-05, 3.3649e-05, 3.4737e-05, 3.5702e-05, 3.6374e-05, 3.6764e-05, 
    3.6796e-05, 3.6673e-05, 3.6283e-05, 3.5788e-05, 3.5198e-05, 3.4556e-05, 
    3.3922e-05, 3.3194e-05, 3.2445e-05, 3.1817e-05, 3.1108e-05, 3.0428e-05, 
    2.9835e-05, 2.9284e-05, 2.8817e-05, 2.8418e-05, 2.8106e-05, 2.7949e-05, 
    2.7902e-05, 2.8066e-05, 2.8281e-05, 2.8672e-05, 2.9049e-05, 2.952e-05, 
    2.9948e-05, 3.0353e-05, 3.0696e-05, 3.0999e-05, 3.1282e-05, 3.1679e-05, 
    3.2068e-05, 3.2512e-05, 3.2968e-05, 3.3406e-05, 3.3789e-05, 3.4134e-05, 
    3.4446e-05, 3.4656e-05, 3.4853e-05, 3.4856e-05, 3.4763e-05, 3.4448e-05, 
    3.4038e-05, 3.3548e-05, 3.2951e-05, 3.2183e-05, 3.142e-05, 3.0496e-05, 
    2.9404e-05, 2.8292e-05, 2.7018e-05, 2.5669e-05, 2.419e-05, 2.2708e-05, 
    2.1143e-05, 1.9683e-05, 1.8377e-05, 1.7323e-05, 1.6597e-05, 1.5993e-05, 
    1.5461e-05, 1.5022e-05, 1.4734e-05, 1.4458e-05, 1.4301e-05, 1.4292e-05, 
    1.4409e-05, 1.4724e-05, 1.517e-05, 1.5717e-05, 1.642e-05, 1.7155e-05, 
    1.7915e-05, 1.8706e-05, 1.9452e-05, 2.0151e-05, 2.0689e-05, 2.1031e-05, 
    2.1171e-05, 2.1121e-05, 2.1049e-05, 2.1001e-05, 2.1029e-05, 2.1258e-05, 
    2.1573e-05, 2.1871e-05, 2.2049e-05, 2.1968e-05, 2.1682e-05, 2.1197e-05, 
    2.0653e-05, 2.0006e-05, 1.9415e-05, 1.8933e-05, 1.8548e-05, 1.8329e-05, 
    1.812e-05, 1.7897e-05, 1.7734e-05, 1.7598e-05, 1.7539e-05, 1.7648e-05, 
    1.7771e-05, 1.796e-05, 1.8217e-05, 1.8519e-05, 1.8791e-05, 1.9269e-05, 
    1.9843e-05, 2.0573e-05, 2.1452e-05, 2.2421e-05, 2.3548e-05, 2.4728e-05, 
    2.6067e-05, 2.7366e-05, 2.874e-05, 3.0105e-05, 3.1465e-05, 3.29e-05, 
    3.4361e-05, 3.5775e-05, 3.7158e-05, 3.8537e-05, 3.9905e-05, 4.1223e-05, 
    4.2516e-05, 4.3704e-05, 4.4729e-05, 4.5639e-05, 4.6336e-05, 4.6879e-05, 
    4.7281e-05, 4.7518e-05, 4.7593e-05, 4.7547e-05, 4.7325e-05, 4.6855e-05, 
    4.6088e-05, 4.4883e-05, 4.3275e-05, 4.1391e-05, 3.9404e-05, 3.736e-05, 
    3.5452e-05, 3.3671e-05, 3.1978e-05, 3.0334e-05, 2.8773e-05, 2.7353e-05, 
    2.6141e-05, 2.5175e-05, 2.4387e-05, 2.3733e-05, 2.3112e-05, 2.2535e-05, 
    2.2016e-05, 2.1531e-05, 2.0985e-05, 2.0475e-05, 1.9926e-05, 1.9483e-05, 
    1.92e-05, 1.9083e-05, 1.913e-05, 1.9401e-05, 1.9851e-05, 2.0464e-05, 
    2.1278e-05, 2.2104e-05, 2.3081e-05, 2.4052e-05, 2.4982e-05, 2.6029e-05, 
    2.6974e-05, 2.7969e-05, 2.8929e-05, 2.9944e-05, 3.0853e-05, 3.1659e-05, 
    3.228e-05, 3.268e-05, 3.2897e-05, 3.2827e-05, 3.2441e-05, 3.183e-05, 
    3.0994e-05, 2.9966e-05, 2.871e-05, 2.7323e-05, 2.5789e-05, 2.4182e-05, 
    2.2485e-05, 2.0819e-05, 1.9204e-05, 1.7655e-05, 1.6237e-05, 1.5083e-05, 
    1.4131e-05, 1.3391e-05, 1.2777e-05, 1.2217e-05, 1.1706e-05, 1.1286e-05, 
    1.0976e-05, 1.0811e-05, 1.0749e-05, 1.0696e-05, 1.0659e-05, 1.0632e-05, 
    1.0623e-05, 1.0699e-05, 1.1167e-05, 1.1882e-05, 1.2935e-05, 1.4191e-05, 
    1.5496e-05, 1.6796e-05, 1.806e-05, 1.9239e-05, 2.035e-05, 2.1398e-05, 
    2.2367e-05, 2.3179e-05, 2.3869e-05, 2.4487e-05, 2.4998e-05, 2.5343e-05, 
    2.578e-05, 2.6221e-05, 2.666e-05, 2.7175e-05, 2.7767e-05, 2.8352e-05, 
    2.9059e-05, 2.9694e-05, 3.0329e-05, 3.0946e-05, 3.1601e-05, 3.2221e-05, 
    3.283e-05, 3.3451e-05, 3.4057e-05, 3.4669e-05, 3.5271e-05, 3.5875e-05, 
    3.6482e-05, 3.7051e-05, 3.7447e-05, 3.7632e-05, 3.767e-05, 3.7522e-05, 
    3.7257e-05, 3.6777e-05, 3.618e-05, 3.5533e-05, 3.468e-05, 3.3639e-05, 
    3.2457e-05, 3.1083e-05, 2.9624e-05, 2.8129e-05, 2.6525e-05, 2.4806e-05, 
    2.3083e-05, 2.1415e-05, 1.9843e-05, 1.8299e-05, 1.6954e-05, 1.5866e-05, 
    1.4964e-05, 1.4297e-05, 1.369e-05, 1.349e-05, 1.3536e-05, 1.3907e-05, 
    1.4544e-05, 1.5346e-05, 1.6452e-05, 1.7745e-05, 1.9114e-05, 2.0567e-05, 
    2.2105e-05, 2.3684e-05, 2.5172e-05, 2.6494e-05, 2.7734e-05, 2.875e-05, 
    2.946e-05, 2.9909e-05, 3.0078e-05, 3.0083e-05, 2.9907e-05, 2.9613e-05, 
    2.909e-05, 2.8438e-05, 2.7654e-05, 2.6812e-05, 2.593e-05, 2.5031e-05, 
    2.4085e-05, 2.3127e-05, 2.228e-05, 2.1369e-05, 2.0493e-05, 1.9716e-05, 
    1.8993e-05, 1.8451e-05, 1.8136e-05, 1.7853e-05, 1.7667e-05, 1.7661e-05, 
    1.7646e-05, 1.7709e-05, 1.7848e-05, 1.8011e-05, 1.8413e-05, 1.8977e-05, 
    1.9532e-05, 2.0175e-05, 2.0808e-05, 2.1463e-05, 2.2142e-05, 2.2788e-05, 
    2.3225e-05, 2.3652e-05, 2.3996e-05, 2.4219e-05, 2.4229e-05, 2.4087e-05, 
    2.3853e-05, 2.353e-05, 2.3129e-05, 2.2572e-05, 2.2009e-05, 2.1435e-05, 
    2.087e-05, 2.0283e-05, 1.9638e-05, 1.9077e-05, 1.8625e-05, 1.8144e-05, 
    1.785e-05, 1.7616e-05, 1.7586e-05, 1.7659e-05, 1.7842e-05, 1.8174e-05, 
    1.8483e-05, 1.8909e-05, 1.924e-05, 1.9573e-05, 1.9939e-05, 2.0378e-05, 
    2.0911e-05, 2.1334e-05, 2.1716e-05, 2.1998e-05, 2.2265e-05, 2.2542e-05, 
    2.2769e-05, 2.2929e-05, 2.3017e-05, 2.3207e-05, 2.3226e-05, 2.3256e-05, 
    2.3256e-05, 2.3177e-05, 2.3082e-05, 2.2955e-05, 2.282e-05, 2.2647e-05, 
    2.26e-05, 2.2512e-05, 2.2557e-05, 2.2634e-05, 2.2798e-05, 2.3013e-05, 
    2.336e-05, 2.3691e-05, 2.4098e-05, 2.4464e-05, 2.4901e-05, 2.5369e-05, 
    2.5948e-05, 2.6463e-05, 2.7125e-05, 2.7758e-05, 2.8401e-05, 2.905e-05, 
    2.9736e-05, 3.0414e-05, 3.1049e-05, 3.1682e-05, 3.2142e-05, 3.2444e-05, 
    3.2494e-05, 3.242e-05, 3.21e-05, 3.1653e-05, 3.1088e-05, 3.0342e-05, 
    2.9453e-05, 2.8632e-05, 2.7743e-05, 2.6853e-05, 2.6081e-05, 2.5398e-05, 
    2.4775e-05, 2.4173e-05, 2.3787e-05, 2.3466e-05, 2.3376e-05, 2.3483e-05, 
    2.3819e-05, 2.448e-05, 2.5281e-05, 2.6212e-05, 2.7254e-05, 2.837e-05, 
    2.9596e-05, 3.0672e-05, 3.1722e-05, 3.2625e-05, 3.3383e-05, 3.393e-05, 
    3.4306e-05, 3.4451e-05, 3.4356e-05, 3.406e-05, 3.3507e-05, 3.2785e-05, 
    3.1836e-05, 3.0702e-05, 2.9513e-05, 2.8288e-05, 2.693e-05, 2.5533e-05, 
    2.4001e-05, 2.2408e-05, 2.0859e-05, 1.9308e-05, 1.7642e-05, 1.6119e-05, 
    1.4511e-05, 1.3045e-05, 1.1625e-05, 1.0251e-05, 8.938e-06, 7.753e-06, 
    6.694e-06, 5.918e-06, 5.485e-06, 5.416e-06, 5.765e-06, 6.442e-06, 
    7.534e-06, 8.816e-06, 1.0323e-05, 1.213e-05, 1.4087e-05, 1.6107e-05, 
    1.8183e-05, 2.0224e-05, 2.2078e-05, 2.3812e-05, 2.5395e-05, 2.6836e-05, 
    2.8092e-05, 2.9072e-05, 2.9865e-05, 3.0368e-05, 3.0376e-05, 3.0093e-05, 
    2.9425e-05, 2.8389e-05, 2.7167e-05, 2.5807e-05, 2.4366e-05, 2.288e-05, 
    2.1317e-05, 1.9915e-05, 1.8496e-05,
  0.022189, 0.02217, 0.022151, 0.02213, 0.022112, 0.022093, 0.022075, 
    0.022057, 0.022038, 0.022019, 0.022001, 0.021982, 0.021963, 0.021943, 
    0.021921, 0.021901, 0.02188, 0.021858, 0.021834, 0.021811, 0.021787, 
    0.021764, 0.021742, 0.021721, 0.021699, 0.021677, 0.021656, 0.021633, 
    0.021609, 0.021586, 0.021564, 0.021544, 0.021525, 0.021508, 0.021492, 
    0.021478, 0.021466, 0.021454, 0.021441, 0.021427, 0.021415, 0.021403, 
    0.021393, 0.021383, 0.021375, 0.021369, 0.021364, 0.021358, 0.021352, 
    0.021346, 0.02134, 0.021334, 0.021329, 0.021324, 0.021318, 0.021312, 
    0.021305, 0.021297, 0.021288, 0.021278, 0.021269, 0.021259, 0.021249, 
    0.021237, 0.021224, 0.02121, 0.021195, 0.021178, 0.021158, 0.021142, 
    0.021124, 0.021105, 0.021087, 0.021069, 0.021051, 0.021033, 0.021017, 
    0.021, 0.020983, 0.020965, 0.020948, 0.020931, 0.020913, 0.020897, 
    0.020882, 0.020863, 0.020845, 0.020827, 0.020808, 0.020791, 0.020769, 
    0.020749, 0.020729, 0.020709, 0.020688, 0.020674, 0.020659, 0.020647, 
    0.020636, 0.020621, 0.02061, 0.020598, 0.020587, 0.020577, 0.020568, 
    0.020557, 0.020553, 0.020547, 0.020541, 0.020535, 0.020524, 0.020517, 
    0.02051, 0.020504, 0.020498, 0.020491, 0.020484, 0.020476, 0.020468, 
    0.020461, 0.020449, 0.020437, 0.020425, 0.020413, 0.020399, 0.020385, 
    0.02037, 0.020355, 0.020339, 0.020319, 0.020301, 0.020282, 0.02026, 
    0.020235, 0.020209, 0.020181, 0.020153, 0.020123, 0.020093, 0.020062, 
    0.020031, 0.019998, 0.019967, 0.019936, 0.019908, 0.01988, 0.019851, 
    0.019822, 0.019791, 0.01976, 0.019734, 0.019706, 0.019679, 0.019652, 
    0.019623, 0.019593, 0.019568, 0.019544, 0.01952, 0.019498, 0.019471, 
    0.019447, 0.019421, 0.019395, 0.019369, 0.019342, 0.019312, 0.019285, 
    0.019257, 0.019229, 0.019201, 0.01917, 0.019143, 0.019117, 0.019091, 
    0.019065, 0.01904, 0.019015, 0.018991, 0.018966, 0.018947, 0.018925, 
    0.018903, 0.018883, 0.018863, 0.018844, 0.018828, 0.018809, 0.018794, 
    0.018783, 0.018775, 0.018768, 0.018762, 0.018755, 0.018752, 0.018751, 
    0.018748, 0.018746, 0.018745, 0.018746, 0.018746, 0.018748, 0.018744, 
    0.018742, 0.01874, 0.018736, 0.018732, 0.018728, 0.018725, 0.01872, 
    0.018711, 0.018701, 0.018692, 0.018683, 0.018672, 0.018658, 0.018645, 
    0.018626, 0.018609, 0.018591, 0.018575, 0.018559, 0.018541, 0.018522, 
    0.018501, 0.018479, 0.018454, 0.018434, 0.018412, 0.018385, 0.018357, 
    0.018327, 0.018296, 0.018265, 0.018238, 0.01821, 0.01818, 0.01815, 
    0.018119, 0.018087, 0.018055, 0.018027, 0.018001, 0.017975, 0.017949, 
    0.017923, 0.017897, 0.017873, 0.017845, 0.017815, 0.017787, 0.017761, 
    0.017735, 0.017712, 0.017685, 0.017663, 0.017641, 0.017617, 0.017595, 
    0.017576, 0.017561, 0.017546, 0.017534, 0.017518, 0.017505, 0.017493, 
    0.017478, 0.01746, 0.017441, 0.017422, 0.017402, 0.017379, 0.017357, 
    0.017335, 0.017314, 0.017294, 0.017274, 0.017256, 0.017233, 0.017211, 
    0.01719, 0.017171, 0.017156, 0.017142, 0.017129, 0.017116, 0.017103, 
    0.017088, 0.017078, 0.01707, 0.017058, 0.017046, 0.017035, 0.017025, 
    0.017012, 0.017006, 0.016999, 0.016991, 0.016981, 0.016967, 0.016949, 
    0.016928, 0.016907, 0.016884, 0.016861, 0.016836, 0.01681, 0.016784, 
    0.016761, 0.016737, 0.016709, 0.016683, 0.01666, 0.016635, 0.01661, 
    0.016583, 0.016557, 0.016528, 0.016497, 0.016465, 0.016434, 0.016404, 
    0.016375, 0.016346, 0.016318, 0.016291, 0.016269, 0.016249, 0.016231, 
    0.016215, 0.016201, 0.016189, 0.016178, 0.016169, 0.016161, 0.016153, 
    0.016146, 0.016139, 0.016132, 0.016123, 0.016114, 0.016104, 0.016092, 
    0.016081, 0.016071, 0.016061, 0.016048, 0.016032, 0.016015, 0.015996, 
    0.015977, 0.01596, 0.01594, 0.015918, 0.015895, 0.015871, 0.015848, 
    0.015826, 0.015803, 0.01578, 0.015756, 0.015731, 0.015707, 0.015683, 
    0.015659, 0.015634, 0.015607, 0.015578, 0.015546, 0.01552, 0.015493, 
    0.015461, 0.01543, 0.015405, 0.015382, 0.01536, 0.015338, 0.015318, 
    0.015301, 0.015283, 0.015265, 0.015249, 0.015232, 0.015217, 0.015201, 
    0.015188, 0.015176, 0.015164, 0.015151, 0.015135, 0.015121, 0.015108, 
    0.015096, 0.015081, 0.015072, 0.015063, 0.015056, 0.015046, 0.015037, 
    0.015029, 0.015022, 0.015013, 0.015007, 0.015002, 0.014998, 0.014991, 
    0.014987, 0.014982, 0.014974, 0.014964, 0.014948, 0.014932, 0.014918, 
    0.014903, 0.014886, 0.014868, 0.01485, 0.014831, 0.014812, 0.014789, 
    0.014765, 0.014739, 0.014712, 0.014682, 0.014653, 0.014623, 0.014596, 
    0.014565, 0.014532, 0.014495, 0.014464, 0.01443, 0.014396, 0.014359, 
    0.014325, 0.014293, 0.014263, 0.014235, 0.011673, 0.011652, 0.011632, 
    0.011613, 0.011593, 0.011575, 0.011552, 0.011538, 0.011516, 0.011496, 
    0.011476, 0.011457, 0.011434, 0.011414, 0.011395, 0.011374, 0.01135, 
    0.011328, 0.01131, 0.011284, 0.011259, 0.011234, 0.01121, 0.011188, 
    0.011165, 0.011144, 0.011123, 0.011103, 0.011085, 0.011066, 0.011048, 
    0.011031, 0.011018, 0.011003, 0.010989, 0.010973, 0.01096, 0.010948, 
    0.010936, 0.010923, 0.010912, 0.010902, 0.010893, 0.010884, 0.010876, 
    0.010864, 0.010856, 0.010848, 0.01084, 0.010832, 0.010826, 0.010818, 
    0.010805, 0.010791, 0.010779, 0.010768, 0.010757, 0.010745, 0.010733, 
    0.010719, 0.010705, 0.010689, 0.010673, 0.010656, 0.010638, 0.010621, 
    0.010604, 0.010582, 0.010566, 0.010547, 0.010528, 0.01051, 0.010492, 
    0.010474, 0.010456, 0.010439, 0.010422, 0.010405, 0.010388, 0.010377, 
    0.01036, 0.010343, 0.010325, 0.010308, 0.010291, 0.010274, 0.010258, 
    0.010242, 0.010226, 0.01021, 0.010194, 0.010178, 0.010162, 0.010147, 
    0.010133, 0.010119, 0.010106, 0.010092, 0.010078, 0.010064, 0.010049, 
    0.010035, 0.010021, 0.010007, 0.0099935, 0.0099806, 0.0099633, 0.0099479, 
    0.0099327, 0.0099184, 0.0099037, 0.0098904, 0.0098761, 0.0098624, 
    0.0098479, 0.0098332, 0.0098184, 0.009804, 0.0097898, 0.009776, 
    0.0097618, 0.0097473, 0.0097326, 0.0097172, 0.0097021, 0.0096864, 
    0.0096709, 0.0096551, 0.009639, 0.009623, 0.009607, 0.0095912, 0.0095755, 
    0.00956, 0.0095445, 0.0095288, 0.0095129, 0.0094969, 0.0094807, 
    0.0094649, 0.0094491, 0.0094339, 0.0094188, 0.0094044, 0.0093905, 
    0.0093767, 0.0093633, 0.0093495, 0.0093354, 0.0093207, 0.0093058, 
    0.0092902, 0.0092742, 0.0092582, 0.0092421, 0.0092265, 0.0092109, 
    0.0091953, 0.0091797, 0.0091641, 0.0091487, 0.0091333, 0.0091182, 
    0.0091034, 0.009089, 0.0090747, 0.0090606, 0.0090464, 0.0090328, 
    0.0090191, 0.0090064, 0.0089935, 0.0089813, 0.0089684, 0.0089561, 
    0.0089433, 0.0089302, 0.0089169, 0.0089036, 0.0088903, 0.0088771, 
    0.0088627, 0.0088483, 0.0088334, 0.0088182, 0.0088037, 0.0087887, 
    0.0087748, 0.0087607, 0.0087472, 0.008734, 0.0087206, 0.0087075, 
    0.0086945, 0.0086818, 0.0086689, 0.0086559, 0.0086424, 0.0086286, 
    0.008614, 0.0085988, 0.008583, 0.0085664, 0.0085496, 0.0085327, 
    0.0085164, 0.0085003, 0.0084845, 0.0084687, 0.0084527, 0.0084367, 
    0.0084206, 0.0084044, 0.0083881, 0.0083717, 0.0083551, 0.0083384, 
    0.0083216, 0.0083048, 0.0082878, 0.0082711, 0.0082541, 0.008237, 0.00822, 
    0.0082032, 0.0081863, 0.0081695, 0.0081527, 0.0081357, 0.008119, 
    0.0081023, 0.0080857, 0.0080698, 0.0080541, 0.0080389, 0.0080241, 
    0.0080099, 0.0079959, 0.0079823, 0.0079691, 0.0079565, 0.0079446, 
    0.0079316, 0.0079189, 0.0079054, 0.0078913, 0.0078772, 0.0078623, 
    0.0078477, 0.007833, 0.0078182, 0.0078038, 0.0077896, 0.0077755, 
    0.0077617, 0.0077479, 0.0077344, 0.0077212, 0.0077082, 0.0076955, 
    0.007683, 0.0076707, 0.0076585, 0.0076465, 0.0076348, 0.0076233, 
    0.007612, 0.0076008, 0.00759, 0.0075791, 0.0075683, 0.0075574, 0.0075465, 
    0.0075358, 0.0075249, 0.0075141, 0.0075031, 0.0074922, 0.0074809, 
    0.0074694, 0.0074578, 0.0074458, 0.0074333, 0.0074206, 0.0074078, 
    0.0073949, 0.0073817, 0.0073683, 0.0073546, 0.0073404, 0.0073261, 
    0.0073113, 0.0072962, 0.0072811, 0.0072657, 0.0072504, 0.0072353, 
    0.0072201, 0.0072049, 0.0071899, 0.0071749, 0.0071601, 0.0071453, 
    0.0071306, 0.0071162, 0.0071019, 0.0070876, 0.0070734, 0.0070593, 
    0.0070453, 0.0070314, 0.0070176, 0.0070038, 0.0069901, 0.0069766, 
    0.0069629, 0.0069491, 0.0069355, 0.0069219, 0.0069084, 0.0068948, 
    0.0068813, 0.0068677, 0.006854, 0.0068404, 0.0068267, 0.0068131, 
    0.0067995, 0.0067859, 0.0067726, 0.006759, 0.0067455, 0.006732, 
    0.0067185, 0.0067051, 0.0066917, 0.0066784, 0.0066652, 0.0066522, 
    0.0066394, 0.0066266, 0.0066141, 0.0066015, 0.006589, 0.0065768, 
    0.0065646, 0.0065526, 0.0065406, 0.0065287, 0.006517, 0.0065052, 
    0.0064935, 0.0064818, 0.0064699, 0.0064577, 0.0064452, 0.0064326, 
    0.0064198, 0.0064068, 0.0063933, 0.0063798, 0.0063663, 0.0063527, 
    0.0063391, 0.0063254, 0.0063118, 0.0062983, 0.0062847, 0.0062709, 
    0.0062571, 0.0062433, 0.0062297, 0.0062161, 0.0062028, 0.00619, 
    0.0061776, 0.0061659, 0.0061547, 0.0061439, 0.0061336, 0.0061237, 
    0.0061141, 0.0061049, 0.006096, 0.0060872, 0.0060788, 0.0060704, 
    0.0060624, 0.0060544, 0.0060467, 0.0060392, 0.0060315, 0.0060238, 
    0.0060158, 0.0060078, 0.0059994, 0.0059909, 0.0059821, 0.005973, 
    0.0059639, 0.0059546, 0.0059448, 0.0059347, 0.0059242, 0.0059132, 
    0.0059018, 0.00589, 0.0058778, 0.0058654, 0.0058526, 0.0058395, 
    0.0058261, 0.0058125, 0.0057986, 0.0057844, 0.0057699, 0.0057552, 
    0.0057405, 0.0057255, 0.0057103, 0.005695, 0.0056797, 0.0056645, 
    0.0056494, 0.0056343, 0.0056194, 0.0056046, 0.00559, 0.0055753, 
    0.0055606, 0.0055458, 0.0055309, 0.0055158, 0.0055004, 0.0054846, 
    0.0054687, 0.0054528, 0.0054368, 0.0054208, 0.0054048, 0.0053888, 
    0.0053728, 0.0053569, 0.005341, 0.0053254, 0.0053099, 0.0052944, 
    0.005279, 0.0052636, 0.0052484, 0.0052333, 0.0052183, 0.0052034, 
    0.0051886, 0.0051738, 0.005159, 0.0051442, 0.0051293, 0.0051143, 
    0.0050992, 0.0050839, 0.0050687, 0.0050534, 0.005038, 0.0050226, 
    0.0050071, 0.0049914, 0.0049758, 0.0049602, 0.0049447, 0.0049292, 
    0.0049136, 0.0048978, 0.0048817, 0.0048655, 0.004849, 0.0048323, 
    0.0048155, 0.0047987, 0.0047818, 0.0047649, 0.004748, 0.0047314, 
    0.0047149, 0.0046986, 0.0046825, 0.0046666, 0.0046506, 0.0046351, 
    0.0046202, 0.0046054, 0.0045912, 0.0045772, 0.0045633, 0.0045497, 
    0.0045362, 0.004523, 0.00451, 0.0044972, 0.0044843, 0.0044714, 0.0044583, 
    0.004445, 0.0044315, 0.0044176, 0.0044038, 0.0043898, 0.0043756, 
    0.0043612, 0.0043465, 0.0043315, 0.0043165, 0.0043013, 0.0042859, 
    0.0042704, 0.0042549, 0.0042392, 0.0042236, 0.0042081, 0.0041926, 
    0.0041769, 0.0041611, 0.0041453, 0.0041292, 0.0041132, 0.0040972, 
    0.0040813, 0.0040654, 0.0040499, 0.0040347, 0.00402, 0.0040059, 
    0.0039921, 0.0039787, 0.0039655, 0.0039527, 0.0039399, 0.0039273, 
    0.0039148, 0.0039021, 0.0038894, 0.0038768, 0.0038642, 0.0038517, 
    0.0038392, 0.0038268, 0.0038144, 0.0038019, 0.0037891, 0.0037761, 
    0.0037632, 0.0037501, 0.0037372, 0.0037241, 0.0037109, 0.0036977, 
    0.0036845, 0.0036713, 0.0036582, 0.0036453, 0.0036323, 0.0036192, 
    0.0036062, 0.003593, 0.0035799, 0.0035666, 0.0035534, 0.0035403, 
    0.0035273, 0.0035143, 0.0035012, 0.0034881, 0.0034751, 0.0034621, 
    0.0034492, 0.0034364, 0.0034235, 0.0034108, 0.0033982, 0.0033857, 
    0.0033734, 0.0033611, 0.0033487, 0.0033361, 0.0033233, 0.0033105, 
    0.0032976, 0.0032846, 0.0032714, 0.0032579, 0.0032445, 0.003231, 
    0.0032177, 0.0032044, 0.0031911, 0.0031779, 0.0031648, 0.0031516, 
    0.0031386, 0.0031255, 0.0031125, 0.0030995, 0.0030865, 0.0030736, 
    0.0030605, 0.0030475, 0.0030344, 0.0030213, 0.0030082, 0.0029952, 
    0.0029823, 0.0029695, 0.0029568, 0.0029441, 0.0029318, 0.0029195, 
    0.0029074, 0.0028957, 0.0028842, 0.0028731, 0.0028621, 0.0028513, 
    0.0028406, 0.00283, 0.0028194, 0.0028089, 0.0027984, 0.002788, 0.0027777, 
    0.0027673, 0.002757, 0.0027466, 0.0027362, 0.0027258, 0.0027154, 
    0.0027049, 0.0026945, 0.002684, 0.0026736, 0.0026631, 0.0026527, 
    0.0026423, 0.0026319, 0.0026214, 0.0026108, 0.0025999, 0.002589, 
    0.002578, 0.0025669, 0.0025557, 0.0025443, 0.0025328, 0.0025213, 
    0.0025098, 0.0024982, 0.0024867, 0.0024753, 0.0024638, 0.0024523, 
    0.0024408, 0.0024294, 0.0024178, 0.0024063, 0.0023948, 0.0023834, 
    0.002372, 0.0023606, 0.0023493, 0.002338, 0.0023267, 0.0023153, 0.002304, 
    0.0022926, 0.0022812, 0.0022698, 0.0022585, 0.0022472, 0.002236, 
    0.0022249, 0.002214, 0.0022035, 0.0021931, 0.0021828, 0.0021727, 
    0.0021628, 0.002153, 0.0021432, 0.0021335, 0.0021238, 0.0021143, 
    0.0021047, 0.0020951, 0.0020855, 0.0020759, 0.0020662, 0.0020563, 
    0.0020465, 0.0020366, 0.0020267, 0.0020167, 0.0020066, 0.0019967, 
    0.0019867, 0.0019766, 0.0019663, 0.0019559, 0.0019452, 0.0019345, 
    0.0019234, 0.0019124, 0.0019013, 0.0018901, 0.0018789, 0.0018675, 
    0.0018561, 0.0018445, 0.001833, 0.0018215, 0.0018101, 0.0017987, 
    0.0017876, 0.0017766, 0.0017658, 0.0017552, 0.0017448, 0.0017345, 
    0.0017245, 0.0017146, 0.0017049, 0.0016956, 0.0016864, 0.0016775, 
    0.001669, 0.0016606, 0.0016524, 0.0016445, 0.0016366, 0.0016289, 
    0.0016211, 0.0016133, 0.0016056, 0.0015979, 0.0015902, 0.0015825, 
    0.0015749, 0.0015672, 0.0015597, 0.001552, 0.0015444, 0.0015367, 
    0.0015289, 0.0015211, 0.0015134, 0.0015057, 0.0014979, 0.0014901, 
    0.0014822, 0.0014743, 0.0014664, 0.0014584, 0.0014505, 0.0014425, 
    0.0014347, 0.0014268, 0.0014189, 0.0014111, 0.0014033, 0.0013955, 
    0.0013878, 0.0013802, 0.0013725, 0.001365, 0.0013575, 0.0013501, 
    0.0013426, 0.0013352, 0.0013277, 0.0013203, 0.0013128, 0.0013054, 
    0.0012979, 0.0012904, 0.001283, 0.0012756, 0.0012682, 0.0012607, 
    0.0012532, 0.0012456, 0.0012379, 0.0012301, 0.0012223, 0.0012145, 
    0.0012066, 0.0011988, 0.0011909, 0.001183, 0.0011753, 0.0011675, 
    0.0011597, 0.0011519, 0.0011441, 0.0011363, 0.0011285, 0.0011208, 
    0.0011131, 0.0011055, 0.0010979, 0.0010905, 0.0010832, 0.001076, 
    0.001069, 0.001062, 0.0010553, 0.0010486, 0.0010422, 0.0010358, 
    0.0010296, 0.0010235, 0.0010176, 0.0010118, 0.0010063, 0.001001, 
    0.00099604, 0.00099119, 0.00098647, 0.00098178, 0.00097728, 0.00097282, 
    0.00096826, 0.00096376, 0.00095923, 0.00095477, 0.00095022, 0.00094567, 
    0.00094099, 0.00093625, 0.00093145, 0.00092651, 0.00092144, 0.00091617, 
    0.00091076, 0.00090509, 0.00089923, 0.00089331, 0.0008872, 0.0008809, 
    0.00087444, 0.0008678, 0.00086104, 0.0008541, 0.00084703, 0.0008399, 
    0.0008328, 0.00082571, 0.00081859, 0.00081144, 0.00080423, 0.0007971, 
    0.00079003, 0.00078302, 0.00077601, 0.00076906, 0.0007622, 0.00075544, 
    0.00074887, 0.00074239, 0.00073607, 0.0007299, 0.00072392, 0.00071805, 
    0.00071238, 0.00070698, 0.00070178, 0.0006968, 0.0006919, 0.00068724, 
    0.00068277, 0.00067844, 0.00067413, 0.00066991, 0.00066577, 0.00066172, 
    0.00065775, 0.00065381, 0.00064989, 0.00064593, 0.00064191, 0.00063791, 
    0.00063381, 0.00062965, 0.00062542, 0.00062096, 0.00061649, 0.00061182, 
    0.0006071, 0.00060228, 0.00059738, 0.00059249, 0.00058758, 0.00058278, 
    0.00057806, 0.00057342, 0.00056888, 0.00056434, 0.00055988, 0.00055545, 
    0.00055106, 0.00054671, 0.00054239, 0.00053816, 0.00053403, 0.00052994, 
    0.00052584, 0.00052189, 0.00051813, 0.00051448, 0.00051097, 0.00050752, 
    0.00050419, 0.00050102, 0.00049789, 0.00049481, 0.0004918, 0.00048885, 
    0.00048593, 0.00048299, 0.00047999, 0.00047699, 0.00047396, 0.00047093, 
    0.00046784, 0.00046462, 0.00046138, 0.00045808, 0.00045473, 0.00045119, 
    0.0004476, 0.00044395, 0.00044029, 0.0004366, 0.00043286, 0.00042914, 
    0.00042552, 0.00042188, 0.00041838, 0.0004149, 0.00041148, 0.00040824, 
    0.00040504, 0.00040192, 0.00039891, 0.00039599, 0.00039312, 0.00039031, 
    0.00038753, 0.00038479, 0.00038214, 0.0003796, 0.00037703, 0.00037454, 
    0.00037211, 0.00036973, 0.00036749, 0.00036533, 0.0003632, 0.00036104, 
    0.00035887, 0.00035676, 0.0003547, 0.00035265, 0.00035063, 0.00034876, 
    0.00034692, 0.00034506, 0.0003432, 0.00034137, 0.00033951, 0.00033764, 
    0.00033576, 0.00033395, 0.00033212, 0.00033032, 0.00032851, 0.00032677, 
    0.00032504, 0.00032337, 0.00032166, 0.00031986, 0.00031799, 0.00031601, 
    0.00031401, 0.00031188, 0.00030965, 0.00030731, 0.00030488, 0.00030236, 
    0.00029973, 0.00029698, 0.00029414, 0.00029126, 0.00028831, 0.00028526, 
    0.00028213, 0.00027894, 0.00027567, 0.00027248, 0.00026923, 0.00026598, 
    0.00026285, 0.00025971, 0.00025668, 0.00025368, 0.00025074, 0.00024797, 
    0.00024521, 0.00024256, 0.00023997, 0.00023741, 0.00023507, 0.00023281, 
    0.00023072, 0.0002288, 0.00022699, 0.00022539, 0.00022399, 0.00022266, 
    0.00022132, 0.0002201, 0.00021888, 0.00021772, 0.0002166, 0.00021557, 
    0.00021463, 0.00021376, 0.00021289, 0.00021201, 0.00021109, 0.00021009, 
    0.00020896, 0.00020775, 0.00020647, 0.00020509, 0.00020364, 0.00020214, 
    0.00020061, 0.00019905, 0.00019745, 0.00019584, 0.00019419, 0.00019256, 
    0.00019091, 0.0001893, 0.00018772, 0.00018616, 0.00018461, 0.00018313, 
    0.00018166, 0.00018032, 0.00017909, 0.00017793, 0.00017687, 0.00017584, 
    0.00017488, 0.0001739, 0.00017298, 0.00017212, 0.00017132, 0.00017052, 
    0.00016976, 0.00016896, 0.00016816, 0.0001674, 0.00016661, 0.00016573, 
    0.00016488, 0.0001639, 0.00016291, 0.00016179, 0.00016058, 0.00015936, 
    0.00015803, 0.00015671, 0.00015527, 0.00015378, 0.00015224, 0.00015078, 
    0.00014929, 0.00014773, 0.00014618, 0.00014465, 0.00014308, 0.00014155, 
    0.00014007, 0.00013865, 0.00013731, 0.00013601, 0.00013476, 0.00013356, 
    0.00013239, 0.00013132, 0.00013026, 0.00012929, 0.0001284, 0.0001275, 
    0.00012666, 0.00012591, 0.00012517, 0.00012446, 0.00012375, 0.0001231, 
    0.00012244, 0.00012179, 0.0001211, 0.00012042, 0.00011976, 0.000119, 
    0.00011817, 0.00011725, 0.00011618, 0.00011516, 0.00011404, 0.00011286, 
    0.00011168, 0.00011043, 0.00010912, 0.00010779, 0.0001065, 0.0001052, 
    0.0001039, 0.00010261, 0.00010135, 0.00010011, 9.898e-05, 9.7905e-05, 
    9.6851e-05, 9.5872e-05, 9.4819e-05, 9.3797e-05, 9.2714e-05, 9.1686e-05, 
    9.0734e-05, 8.9782e-05, 8.8917e-05, 8.8053e-05, 8.7292e-05, 8.6581e-05, 
    8.5998e-05, 8.5514e-05, 8.5088e-05, 8.4735e-05, 8.4488e-05, 8.431e-05, 
    8.4283e-05, 8.4276e-05, 8.4461e-05, 8.4737e-05, 8.5147e-05, 8.5627e-05, 
    8.6138e-05, 8.6623e-05, 8.7141e-05, 8.7604e-05, 8.8035e-05, 8.8444e-05, 
    8.8792e-05, 8.9085e-05, 8.9297e-05, 8.9339e-05, 8.9287e-05, 8.9025e-05, 
    8.8758e-05, 8.8383e-05, 8.793e-05, 8.742e-05, 8.6878e-05, 8.6327e-05, 
    8.5737e-05, 8.5147e-05, 8.449e-05, 8.3635e-05, 8.2747e-05, 8.1737e-05, 
    8.0595e-05, 7.9486e-05, 7.8216e-05, 7.6924e-05, 7.5585e-05, 7.4195e-05, 
    7.2882e-05, 7.1453e-05, 7.0007e-05, 6.8624e-05, 6.7241e-05, 6.589e-05, 
    6.4563e-05, 6.3325e-05, 6.2242e-05, 6.1237e-05, 6.0312e-05, 5.9501e-05, 
    5.8714e-05, 5.8023e-05, 5.7403e-05, 5.6811e-05, 5.6186e-05, 5.5597e-05, 
    5.5033e-05, 5.4507e-05, 5.4024e-05, 5.3556e-05, 5.3128e-05, 5.2688e-05, 
    5.2159e-05, 5.1628e-05, 5.1018e-05, 5.0352e-05, 4.9658e-05, 4.9021e-05, 
    4.8402e-05, 4.7876e-05, 4.7351e-05, 4.6856e-05, 4.6384e-05, 4.5952e-05, 
    4.5569e-05, 4.5196e-05, 4.4984e-05, 4.4823e-05, 4.471e-05, 4.4688e-05, 
    4.4645e-05, 4.4635e-05, 4.4635e-05, 4.471e-05, 4.4687e-05, 4.4703e-05, 
    4.4719e-05, 4.4769e-05, 4.4875e-05, 4.4914e-05, 4.4909e-05, 4.4977e-05, 
    4.5037e-05, 4.5053e-05, 4.5148e-05, 4.5174e-05, 4.5199e-05, 4.5288e-05, 
    4.5341e-05, 4.5474e-05, 4.5599e-05, 4.5745e-05, 4.5929e-05, 4.6125e-05, 
    4.6259e-05, 4.6239e-05, 4.615e-05, 4.6047e-05, 4.5999e-05, 4.5968e-05, 
    4.6001e-05, 4.5987e-05, 4.5788e-05, 4.5557e-05, 4.5246e-05, 4.4779e-05, 
    4.4261e-05, 4.3713e-05, 4.3152e-05, 4.2571e-05, 4.2138e-05, 4.1787e-05, 
    4.1546e-05, 4.1401e-05, 4.1361e-05, 4.1433e-05, 4.1621e-05, 4.2035e-05, 
    4.2627e-05, 4.3446e-05, 4.449e-05, 4.575e-05, 4.7139e-05, 4.863e-05, 
    5.0205e-05, 5.1828e-05, 5.3408e-05, 5.4959e-05, 5.6418e-05, 5.7816e-05, 
    5.9098e-05, 6.0245e-05, 6.1169e-05, 6.1863e-05, 6.2457e-05, 6.2785e-05, 
    6.2959e-05, 6.3e-05, 6.2789e-05, 6.2447e-05, 6.1804e-05, 6.0923e-05, 
    5.9836e-05, 5.8535e-05, 5.7021e-05, 5.5294e-05, 5.3332e-05, 5.12e-05, 
    4.9038e-05, 4.6736e-05, 4.4393e-05, 4.1994e-05, 3.9615e-05, 3.7196e-05, 
    3.4868e-05, 3.264e-05, 3.0375e-05, 2.8303e-05, 2.6416e-05, 2.4736e-05, 
    2.3378e-05, 2.2441e-05, 2.1756e-05, 2.1212e-05, 2.0982e-05, 2.0907e-05, 
    2.0943e-05, 2.1208e-05, 2.1578e-05, 2.2065e-05, 2.2664e-05, 2.3445e-05, 
    2.4379e-05, 2.5398e-05, 2.6485e-05, 2.7499e-05, 2.8489e-05, 2.9313e-05, 
    3.0188e-05, 3.0942e-05, 3.1696e-05, 3.2403e-05, 3.3072e-05, 3.366e-05, 
    3.4128e-05, 3.4551e-05, 3.4898e-05, 3.5121e-05, 3.5216e-05, 3.5245e-05, 
    3.5159e-05, 3.4919e-05, 3.4536e-05, 3.3996e-05, 3.3327e-05, 3.255e-05, 
    3.1723e-05, 3.0776e-05, 2.9928e-05, 2.8919e-05, 2.8077e-05, 2.7274e-05, 
    2.6531e-05, 2.5889e-05, 2.5287e-05, 2.4773e-05, 2.4293e-05, 2.3868e-05, 
    2.3358e-05, 2.2963e-05, 2.2622e-05, 2.2363e-05, 2.2192e-05, 2.2102e-05, 
    2.1977e-05, 2.191e-05, 2.1872e-05, 2.1736e-05, 2.17e-05, 2.1769e-05, 
    2.1931e-05, 2.2176e-05, 2.2615e-05, 2.3168e-05, 2.3806e-05, 2.4608e-05, 
    2.5596e-05, 2.6692e-05, 2.789e-05, 2.9077e-05, 3.0257e-05, 3.137e-05, 
    3.2505e-05, 3.3649e-05, 3.4737e-05, 3.5702e-05, 3.6374e-05, 3.6764e-05, 
    3.6796e-05, 3.6673e-05, 3.6283e-05, 3.5788e-05, 3.5198e-05, 3.4556e-05, 
    3.3922e-05, 3.3194e-05, 3.2445e-05, 3.1817e-05, 3.1108e-05, 3.0428e-05, 
    2.9835e-05, 2.9284e-05, 2.8817e-05, 2.8418e-05, 2.8106e-05, 2.7949e-05, 
    2.7902e-05, 2.8066e-05, 2.8281e-05, 2.8672e-05, 2.9049e-05, 2.952e-05, 
    2.9948e-05, 3.0353e-05, 3.0696e-05, 3.0999e-05, 3.1282e-05, 3.1679e-05, 
    3.2068e-05, 3.2512e-05, 3.2968e-05, 3.3406e-05, 3.3789e-05, 3.4134e-05, 
    3.4446e-05, 3.4656e-05, 3.4853e-05, 3.4856e-05, 3.4763e-05, 3.4448e-05, 
    3.4038e-05, 3.3548e-05, 3.2951e-05, 3.2183e-05, 3.142e-05, 3.0496e-05, 
    2.9404e-05, 2.8292e-05, 2.7018e-05, 2.5669e-05, 2.419e-05, 2.2708e-05, 
    2.1143e-05, 1.9683e-05, 1.8377e-05, 1.7323e-05, 1.6597e-05, 1.5993e-05, 
    1.5461e-05, 1.5022e-05, 1.4734e-05, 1.4458e-05, 1.4301e-05, 1.4292e-05, 
    1.4409e-05, 1.4724e-05, 1.517e-05, 1.5717e-05, 1.642e-05, 1.7155e-05, 
    1.7915e-05, 1.8706e-05, 1.9452e-05, 2.0151e-05, 2.0689e-05, 2.1031e-05, 
    2.1171e-05, 2.1121e-05, 2.1049e-05, 2.1001e-05, 2.1029e-05, 2.1258e-05, 
    2.1573e-05, 2.1871e-05, 2.2049e-05, 2.1968e-05, 2.1682e-05, 2.1197e-05, 
    2.0653e-05, 2.0006e-05, 1.9415e-05, 1.8933e-05, 1.8548e-05, 1.8329e-05, 
    1.812e-05, 1.7897e-05, 1.7734e-05, 1.7598e-05, 1.7539e-05, 1.7648e-05, 
    1.7771e-05, 1.796e-05, 1.8217e-05, 1.8519e-05, 1.8791e-05, 1.9269e-05, 
    1.9843e-05, 2.0573e-05, 2.1452e-05, 2.2421e-05, 2.3548e-05, 2.4728e-05, 
    2.6067e-05, 2.7366e-05, 2.874e-05, 3.0105e-05, 3.1465e-05, 3.29e-05, 
    3.4361e-05, 3.5775e-05, 3.7158e-05, 3.8537e-05, 3.9905e-05, 4.1223e-05, 
    4.2516e-05, 4.3704e-05, 4.4729e-05, 4.5639e-05, 4.6336e-05, 4.6879e-05, 
    4.7281e-05, 4.7518e-05, 4.7593e-05, 4.7547e-05, 4.7325e-05, 4.6855e-05, 
    4.6088e-05, 4.4883e-05, 4.3275e-05, 4.1391e-05, 3.9404e-05, 3.736e-05, 
    3.5452e-05, 3.3671e-05, 3.1978e-05, 3.0334e-05, 2.8773e-05, 2.7353e-05, 
    2.6141e-05, 2.5175e-05, 2.4387e-05, 2.3733e-05, 2.3112e-05, 2.2535e-05, 
    2.2016e-05, 2.1531e-05, 2.0985e-05, 2.0475e-05, 1.9926e-05, 1.9483e-05, 
    1.92e-05, 1.9083e-05, 1.913e-05, 1.9401e-05, 1.9851e-05, 2.0464e-05, 
    2.1278e-05, 2.2104e-05, 2.3081e-05, 2.4052e-05, 2.4982e-05, 2.6029e-05, 
    2.6974e-05, 2.7969e-05, 2.8929e-05, 2.9944e-05, 3.0853e-05, 3.1659e-05, 
    3.228e-05, 3.268e-05, 3.2897e-05, 3.2827e-05, 3.2441e-05, 3.183e-05, 
    3.0994e-05, 2.9966e-05, 2.871e-05, 2.7323e-05, 2.5789e-05, 2.4182e-05, 
    2.2485e-05, 2.0819e-05, 1.9204e-05, 1.7655e-05, 1.6237e-05, 1.5083e-05, 
    1.4131e-05, 1.3391e-05, 1.2777e-05, 1.2217e-05, 1.1706e-05, 1.1286e-05, 
    1.0976e-05, 1.0811e-05, 1.0749e-05, 1.0696e-05, 1.0659e-05, 1.0632e-05, 
    1.0623e-05, 1.0699e-05, 1.1167e-05, 1.1882e-05, 1.2935e-05, 1.4191e-05, 
    1.5496e-05, 1.6796e-05, 1.806e-05, 1.9239e-05, 2.035e-05, 2.1398e-05, 
    2.2367e-05, 2.3179e-05, 2.3869e-05, 2.4487e-05, 2.4998e-05, 2.5343e-05, 
    2.578e-05, 2.6221e-05, 2.666e-05, 2.7175e-05, 2.7767e-05, 2.8352e-05, 
    2.9059e-05, 2.9694e-05, 3.0329e-05, 3.0946e-05, 3.1601e-05, 3.2221e-05, 
    3.283e-05, 3.3451e-05, 3.4057e-05, 3.4669e-05, 3.5271e-05, 3.5875e-05, 
    3.6482e-05, 3.7051e-05, 3.7447e-05, 3.7632e-05, 3.767e-05, 3.7522e-05, 
    3.7257e-05, 3.6777e-05, 3.618e-05, 3.5533e-05, 3.468e-05, 3.3639e-05, 
    3.2457e-05, 3.1083e-05, 2.9624e-05, 2.8129e-05, 2.6525e-05, 2.4806e-05, 
    2.3083e-05, 2.1415e-05, 1.9843e-05, 1.8299e-05, 1.6954e-05, 1.5866e-05, 
    1.4964e-05, 1.4297e-05, 1.369e-05, 1.349e-05, 1.3536e-05, 1.3907e-05, 
    1.4544e-05, 1.5346e-05, 1.6452e-05, 1.7745e-05, 1.9114e-05, 2.0567e-05, 
    2.2105e-05, 2.3684e-05, 2.5172e-05, 2.6494e-05, 2.7734e-05, 2.875e-05, 
    2.946e-05, 2.9909e-05, 3.0078e-05, 3.0083e-05, 2.9907e-05, 2.9613e-05, 
    2.909e-05, 2.8438e-05, 2.7654e-05, 2.6812e-05, 2.593e-05, 2.5031e-05, 
    2.4085e-05, 2.3127e-05, 2.228e-05, 2.1369e-05, 2.0493e-05, 1.9716e-05, 
    1.8993e-05, 1.8451e-05, 1.8136e-05, 1.7853e-05, 1.7667e-05, 1.7661e-05, 
    1.7646e-05, 1.7709e-05, 1.7848e-05, 1.8011e-05, 1.8413e-05, 1.8977e-05, 
    1.9532e-05, 2.0175e-05, 2.0808e-05, 2.1463e-05, 2.2142e-05, 2.2788e-05, 
    2.3225e-05, 2.3652e-05, 2.3996e-05, 2.4219e-05, 2.4229e-05, 2.4087e-05, 
    2.3853e-05, 2.353e-05, 2.3129e-05, 2.2572e-05, 2.2009e-05, 2.1435e-05, 
    2.087e-05, 2.0283e-05, 1.9638e-05, 1.9077e-05, 1.8625e-05, 1.8144e-05, 
    1.785e-05, 1.7616e-05, 1.7586e-05, 1.7659e-05, 1.7842e-05, 1.8174e-05, 
    1.8483e-05, 1.8909e-05, 1.924e-05, 1.9573e-05, 1.9939e-05, 2.0378e-05, 
    2.0911e-05, 2.1334e-05, 2.1716e-05, 2.1998e-05, 2.2265e-05, 2.2542e-05, 
    2.2769e-05, 2.2929e-05, 2.3017e-05, 2.3207e-05, 2.3226e-05, 2.3256e-05, 
    2.3256e-05, 2.3177e-05, 2.3082e-05, 2.2955e-05, 2.282e-05, 2.2647e-05, 
    2.26e-05, 2.2512e-05, 2.2557e-05, 2.2634e-05, 2.2798e-05, 2.3013e-05, 
    2.336e-05, 2.3691e-05, 2.4098e-05, 2.4464e-05, 2.4901e-05, 2.5369e-05, 
    2.5948e-05, 2.6463e-05, 2.7125e-05, 2.7758e-05, 2.8401e-05, 2.905e-05, 
    2.9736e-05, 3.0414e-05, 3.1049e-05, 3.1682e-05, 3.2142e-05, 3.2444e-05, 
    3.2494e-05, 3.242e-05, 3.21e-05, 3.1653e-05, 3.1088e-05, 3.0342e-05, 
    2.9453e-05, 2.8632e-05, 2.7743e-05, 2.6853e-05, 2.6081e-05, 2.5398e-05, 
    2.4775e-05, 2.4173e-05, 2.3787e-05, 2.3466e-05, 2.3376e-05, 2.3483e-05, 
    2.3819e-05, 2.448e-05, 2.5281e-05, 2.6212e-05, 2.7254e-05, 2.837e-05, 
    2.9596e-05, 3.0672e-05, 3.1722e-05, 3.2625e-05, 3.3383e-05, 3.393e-05, 
    3.4306e-05, 3.4451e-05, 3.4356e-05, 3.406e-05, 3.3507e-05, 3.2785e-05, 
    3.1836e-05, 3.0702e-05, 2.9513e-05, 2.8288e-05, 2.693e-05, 2.5533e-05, 
    2.4001e-05, 2.2408e-05, 2.0859e-05, 1.9308e-05, 1.7642e-05, 1.6119e-05, 
    1.4511e-05, 1.3045e-05, 1.1625e-05, 1.0251e-05, 8.938e-06, 7.753e-06, 
    6.694e-06, 5.918e-06, 5.485e-06, 5.416e-06, 5.765e-06, 6.442e-06, 
    7.534e-06, 8.816e-06, 1.0323e-05, 1.213e-05, 1.4087e-05, 1.6107e-05, 
    1.8183e-05, 2.0224e-05, 2.2078e-05, 2.3812e-05, 2.5395e-05, 2.6836e-05, 
    2.8092e-05, 2.9072e-05, 2.9865e-05, 3.0368e-05, 3.0376e-05, 3.0093e-05, 
    2.9425e-05, 2.8389e-05, 2.7167e-05, 2.5807e-05, 2.4366e-05, 2.288e-05, 
    2.1317e-05, 1.9915e-05, 1.8496e-05 ;

 bangle_L2 =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 0.002548, 0.0025362, 0.0025243, 
    0.0025124, 0.0025006, 0.0024887, 0.0024771, 0.0024656, 0.0024541, 
    0.0024431, 0.002432, 0.0024207, 0.0024094, 0.0023982, 0.002387, 
    0.0023757, 0.0023646, 0.0023533, 0.0023421, 0.0023309, 0.0023201, 
    0.0023093, 0.0022988, 0.0022881, 0.0022776, 0.0022668, 0.0022561, 
    0.0022454, 0.0022348, 0.0022246, 0.0022149, 0.002205, 0.0021955, 
    0.0021864, 0.0021776, 0.0021688, 0.0021598, 0.0021507, 0.0021414, 
    0.0021324, 0.0021231, 0.0021137, 0.0021044, 0.0020951, 0.002085, 
    0.0020751, 0.0020652, 0.0020548, 0.0020446, 0.002034, 0.0020235, 
    0.0020125, 0.0020016, 0.00199, 0.0019786, 0.0019668, 0.0019546, 
    0.0019426, 0.0019299, 0.0019176, 0.0019048, 0.001892, 0.0018789, 
    0.0018655, 0.001852, 0.0018387, 0.0018254, 0.0018125, 0.0017996, 
    0.0017869, 0.0017745, 0.0017626, 0.001751, 0.0017395, 0.0017287, 
    0.0017185, 0.0017082, 0.0016986, 0.0016895, 0.0016808, 0.0016722, 
    0.0016641, 0.0016563, 0.001649, 0.0016415, 0.0016347, 0.0016279, 
    0.0016212, 0.0016142, 0.0016077, 0.001601, 0.0015947, 0.0015879, 
    0.0015813, 0.0015746, 0.0015681, 0.0015617, 0.001555, 0.001548, 
    0.0015408, 0.0015341, 0.0015269, 0.0015196, 0.0015123, 0.001505, 
    0.0014972, 0.0014901, 0.0014826, 0.0014751, 0.0014678, 0.0014603, 
    0.0014528, 0.0014452, 0.0014376, 0.0014302, 0.0014228, 0.0014151, 
    0.0014076, 0.0014002, 0.0013924, 0.0013846, 0.0013768, 0.0013694, 
    0.0013616, 0.0013537, 0.001346, 0.001338, 0.0013301, 0.0013222, 
    0.0013142, 0.0013063, 0.0012981, 0.0012901, 0.0012818, 0.0012735, 
    0.0012651, 0.0012568, 0.0012483, 0.0012401, 0.001232, 0.0012239, 
    0.0012156, 0.0012076, 0.0011995, 0.0011914, 0.0011831, 0.0011749, 
    0.0011669, 0.0011589, 0.0011509, 0.0011433, 0.0011356, 0.0011279, 
    0.0011205, 0.001113, 0.0011058, 0.0010986, 0.0010916, 0.0010847, 
    0.0010777, 0.0010706, 0.0010642, 0.0010573, 0.0010509, 0.0010447, 
    0.0010385, 0.0010323, 0.0010265, 0.0010209, 0.0010153, 0.0010099, 
    0.0010047, 0.00099967, 0.00099492, 0.00099023, 0.00098577, 0.00098165, 
    0.00097747, 0.00097346, 0.00096921, 0.00096496, 0.00096071, 0.0009564, 
    0.00095231, 0.00094779, 0.00094328, 0.0009388, 0.00093422, 0.00092929, 
    0.00092443, 0.00091934, 0.00091422, 0.00090894, 0.00090347, 0.00089762, 
    0.00089163, 0.00088509, 0.00087858, 0.0008716, 0.00086489, 0.00085803, 
    0.00085102, 0.00084392, 0.00083687, 0.00082974, 0.00082257, 0.0008152, 
    0.00080763, 0.00080024, 0.00079265, 0.00078513, 0.00077787, 0.00077059, 
    0.0007635, 0.0007567, 0.00074981, 0.00074344, 0.00073712, 0.0007311, 
    0.00072531, 0.00071978, 0.00071419, 0.00070906, 0.00070418, 0.0006995, 
    0.00069486, 0.00069081, 0.00068675, 0.0006829, 0.00067922, 0.00067555, 
    0.0006719, 0.00066822, 0.00066453, 0.00066098, 0.00065716, 0.00065331, 
    0.00064953, 0.00064572, 0.00064166, 0.00063712, 0.00063229, 0.00062743, 
    0.00062256, 0.00061757, 0.00061229, 0.00060709, 0.00060163, 0.00059629, 
    0.0005908, 0.00058549, 0.00058026, 0.00057507, 0.00056996, 0.00056498, 
    0.00056028, 0.00055557, 0.00055082, 0.00054615, 0.00054163, 0.00053717, 
    0.00053289, 0.00052852, 0.00052446, 0.00052065, 0.00051692, 0.00051349, 
    0.00051022, 0.00050712, 0.00050424, 0.00050153, 0.00049888, 0.00049618, 
    0.00049333, 0.00049071, 0.00048821, 0.00048562, 0.00048291, 0.00048012, 
    0.00047719, 0.00047399, 0.00047086, 0.00046773, 0.00046458, 0.00046141, 
    0.00045783, 0.00045394, 0.0004503, 0.00044647, 0.00044264, 0.00043889, 
    0.00043517, 0.00043144, 0.00042792, 0.0004245, 0.00042126, 0.00041787, 
    0.00041468, 0.00041159, 0.00040852, 0.00040545, 0.00040245, 0.00039948, 
    0.00039674, 0.00039429, 0.00039192, 0.0003894, 0.00038736, 0.00038523, 
    0.00038307, 0.00038098, 0.00037883, 0.00037665, 0.00037449, 0.00037215, 
    0.00037003, 0.00036803, 0.00036616, 0.00036463, 0.00036301, 0.00036162, 
    0.00036029, 0.00035902, 0.0003578, 0.00035662, 0.00035532, 0.00035394, 
    0.00035249, 0.000351, 0.0003495, 0.00034789, 0.00034628, 0.00034491, 
    0.00034355, 0.00034196, 0.00034038, 0.00033873, 0.00033711, 0.00033538, 
    0.00033371, 0.0003317, 0.00032935, 0.00032688, 0.00032438, 0.00032182, 
    0.00031905, 0.00031606, 0.00031303, 0.00030986, 0.0003064, 0.00030289, 
    0.00029923, 0.00029527, 0.00029133, 0.0002875, 0.00028364, 0.00027992, 
    0.00027622, 0.00027265, 0.00026911, 0.0002658, 0.00026225, 0.0002588, 
    0.00025548, 0.00025222, 0.00024912, 0.00024634, 0.0002436, 0.00024123, 
    0.00023919, 0.00023742, 0.00023573, 0.00023435, 0.00023305, 0.00023188, 
    0.00023072, 0.00022962, 0.00022856, 0.00022752, 0.00022666, 0.00022579, 
    0.00022488, 0.00022413, 0.00022336, 0.00022288, 0.00022234, 0.00022185, 
    0.00022116, 0.00022036, 0.00021949, 0.00021853, 0.00021723, 0.00021562, 
    0.00021411, 0.00021263, 0.00021081, 0.00020896, 0.00020718, 0.00020532, 
    0.00020352, 0.00020196, 0.00020014, 0.00019844, 0.00019676, 0.00019512, 
    0.00019364, 0.00019217, 0.00019085, 0.00018973, 0.0001887, 0.00018772, 
    0.00018687, 0.0001862, 0.00018534, 0.00018464, 0.0001839, 0.00018335, 
    0.00018283, 0.00018235, 0.0001817, 0.000181, 0.00018065, 0.00017997, 
    0.00017915, 0.00017841, 0.00017771, 0.00017679, 0.00017577, 0.00017452, 
    0.0001729, 0.00017133, 0.00016966, 0.00016777, 0.00016597, 0.00016427, 
    0.00016245, 0.00016059, 0.00015877, 0.00015707, 0.00015532, 0.00015359, 
    0.0001518, 0.00015008, 0.00014845, 0.00014673, 0.00014521, 0.00014383, 
    0.00014263, 0.00014139, 0.00014022, 0.0001392, 0.00013844, 0.00013763, 
    0.00013687, 0.00013622, 0.00013565, 0.00013516, 0.00013475, 0.00013424, 
    0.00013373, 0.00013325, 0.00013288, 0.0001322, 0.00013155, 0.00013088, 
    0.00013007, 0.00012929, 0.00012847, 0.0001275, 0.00012645, 0.00012513, 
    0.00012375, 0.00012233, 0.00012076, 0.00011932, 0.0001178, 0.00011578, 
    0.00011418, 0.00011263, 0.00011121, 0.00010966, 0.0001082, 0.00010696, 
    0.0001056, 0.00010405, 0.00010262, 0.00010139, 0.00010028, 9.9289e-05, 
    9.8352e-05, 9.7269e-05, 9.6322e-05, 9.5355e-05, 9.4581e-05, 9.3888e-05, 
    9.3395e-05, 9.2822e-05, 9.2375e-05, 9.215e-05, 9.2274e-05, 9.2429e-05, 
    9.2745e-05, 9.3209e-05, 9.4e-05, 9.4923e-05, 9.5877e-05, 9.6805e-05, 
    9.789e-05, 9.9109e-05, 0.00010036, 0.00010156, 0.00010263, 0.00010375, 
    0.00010442, 0.00010514, 0.00010561, 0.00010587, 0.00010605, 0.00010631, 
    0.00010637, 0.00010625, 0.00010592, 0.00010546, 0.00010479, 0.00010427, 
    0.00010375, 0.00010294, 0.00010221, 0.00010131, 0.00010035, 9.9014e-05, 
    9.7613e-05, 9.5878e-05, 9.4195e-05, 9.2275e-05, 9.0662e-05, 8.895e-05, 
    8.6734e-05, 8.4683e-05, 8.26e-05, 8.0543e-05, 7.855e-05, 7.6785e-05, 
    7.5073e-05, 7.3427e-05, 7.1873e-05, 7.0415e-05, 6.8886e-05, 6.7577e-05, 
    6.6443e-05, 6.5413e-05, 6.4427e-05, 6.3657e-05, 6.2924e-05, 6.2247e-05, 
    6.1582e-05, 6.1078e-05, 6.0515e-05, 5.9845e-05, 5.9185e-05, 5.8599e-05, 
    5.779e-05, 5.7125e-05, 5.6364e-05, 5.5719e-05, 5.5069e-05, 5.4394e-05, 
    5.3517e-05, 5.2559e-05, 5.1677e-05, 5.0936e-05, 5.0524e-05, 5.012e-05, 
    4.9927e-05, 4.9543e-05, 4.9397e-05, 4.9436e-05, 4.9263e-05, 4.9199e-05, 
    4.9321e-05, 4.9631e-05, 4.9917e-05, 5.0107e-05, 5.0077e-05, 5.0002e-05, 
    5.0148e-05, 5.0411e-05, 5.0464e-05, 5.0892e-05, 5.1089e-05, 5.1535e-05, 
    5.1743e-05, 5.222e-05, 5.2405e-05, 5.2622e-05, 5.2804e-05, 5.3277e-05, 
    5.3783e-05, 5.4235e-05, 5.4696e-05, 5.5105e-05, 5.5316e-05, 5.551e-05, 
    5.5772e-05, 5.5965e-05, 5.6215e-05, 5.6583e-05, 5.6922e-05, 5.6966e-05, 
    5.6919e-05, 5.6883e-05, 5.6578e-05, 5.6111e-05, 5.5599e-05, 5.4976e-05, 
    5.4225e-05, 5.3386e-05, 5.2707e-05, 5.2233e-05, 5.1704e-05, 5.1392e-05, 
    5.1276e-05, 5.1244e-05, 5.1634e-05, 5.2083e-05, 5.2729e-05, 5.3195e-05, 
    5.4194e-05, 5.5603e-05, 5.7075e-05, 5.8722e-05, 6.061e-05, 6.2878e-05, 
    6.5221e-05, 6.7812e-05, 7.0325e-05, 7.2923e-05, 7.5713e-05, 7.8212e-05, 
    8.0591e-05, 8.2984e-05, 8.4986e-05, 8.6869e-05, 8.8362e-05, 8.9439e-05, 
    9.0055e-05, 9.0312e-05, 9.0199e-05, 8.9608e-05, 8.8774e-05, 8.7384e-05, 
    8.5764e-05, 8.376e-05, 8.1353e-05, 7.858e-05, 7.5539e-05, 7.2238e-05, 
    6.8849e-05, 6.5368e-05, 6.178e-05, 5.8019e-05, 5.4237e-05, 5.0365e-05, 
    4.6464e-05, 4.2652e-05, 3.9075e-05, 3.5674e-05, 3.2772e-05, 3.0385e-05, 
    2.8111e-05, 2.6242e-05, 2.4846e-05, 2.3637e-05, 2.2767e-05, 2.244e-05, 
    2.2163e-05, 2.2242e-05, 2.2549e-05, 2.308e-05, 2.3761e-05, 2.4746e-05, 
    2.6e-05, 2.7325e-05, 2.9055e-05, 3.1064e-05, 3.3104e-05, 3.5222e-05, 
    3.6899e-05, 3.8647e-05, 4.0339e-05, 4.1715e-05, 4.3029e-05, 4.4071e-05, 
    4.5131e-05, 4.5894e-05, 4.6569e-05, 4.7012e-05, 4.7246e-05, 4.7269e-05, 
    4.7193e-05, 4.6902e-05, 4.6736e-05, 4.6118e-05, 4.5441e-05, 4.4553e-05, 
    4.3532e-05, 4.2481e-05, 4.1169e-05, 3.9896e-05, 3.8586e-05, 3.731e-05, 
    3.5973e-05, 3.4791e-05, 3.3834e-05, 3.2878e-05, 3.1954e-05, 3.1029e-05, 
    3.0196e-05, 2.935e-05, 2.8771e-05, 2.8273e-05, 2.7869e-05, 2.7455e-05, 
    2.7197e-05, 2.6952e-05, 2.6764e-05, 2.6718e-05, 2.6693e-05, 2.6903e-05, 
    2.7309e-05, 2.7876e-05, 2.8471e-05, 2.9398e-05, 3.0578e-05, 3.1815e-05, 
    3.336e-05, 3.4804e-05, 3.644e-05, 3.8328e-05, 4.0526e-05, 4.273e-05, 
    4.5081e-05, 4.7109e-05, 4.8886e-05, 5.0451e-05, 5.166e-05, 5.2413e-05, 
    5.2758e-05, 5.2847e-05, 5.2737e-05, 5.2246e-05, 5.1466e-05, 5.0629e-05, 
    4.9596e-05, 4.8561e-05, 4.7453e-05, 4.6371e-05, 4.5223e-05, 4.4252e-05, 
    4.3123e-05, 4.1988e-05, 4.1053e-05, 4.034e-05, 3.9921e-05, 3.9544e-05, 
    3.9698e-05, 3.9895e-05, 4.0319e-05, 4.0806e-05, 4.1462e-05, 4.228e-05, 
    4.3146e-05, 4.3931e-05, 4.4797e-05, 4.5575e-05, 4.6466e-05, 4.7333e-05, 
    4.8102e-05, 4.8801e-05, 4.9353e-05, 4.9964e-05, 5.057e-05, 5.1119e-05, 
    5.1545e-05, 5.1936e-05, 5.2105e-05, 5.2046e-05, 5.178e-05, 5.1311e-05, 
    5.077e-05, 5.0173e-05, 4.9453e-05, 4.8351e-05, 4.7072e-05, 4.5809e-05, 
    4.4298e-05, 4.2453e-05, 4.0055e-05, 3.7445e-05, 3.459e-05, 3.1961e-05, 
    2.9494e-05, 2.7145e-05, 2.4905e-05, 2.322e-05, 2.1831e-05, 2.0849e-05, 
    2.0119e-05, 1.9498e-05, 1.9124e-05, 1.8659e-05, 1.8586e-05, 1.8453e-05, 
    1.8694e-05, 1.9119e-05, 1.9632e-05, 2.0372e-05, 2.1282e-05, 2.2291e-05, 
    2.3645e-05, 2.4927e-05, 2.6117e-05, 2.7361e-05, 2.8138e-05, 2.8941e-05, 
    2.931e-05, 2.9892e-05, 3.0269e-05, 3.0473e-05, 3.0995e-05, 3.1212e-05, 
    3.1405e-05, 3.1492e-05, 3.138e-05, 3.1295e-05, 3.0839e-05, 3.0424e-05, 
    2.9853e-05, 2.9283e-05, 2.8562e-05, 2.7923e-05, 2.7319e-05, 2.7004e-05, 
    2.6725e-05, 2.647e-05, 2.6549e-05, 2.6697e-05, 2.6838e-05, 2.7158e-05, 
    2.7204e-05, 2.7112e-05, 2.7352e-05, 2.757e-05, 2.7867e-05, 2.8216e-05, 
    2.8964e-05, 2.9958e-05, 3.1267e-05, 3.2757e-05, 3.455e-05, 3.6442e-05, 
    3.8544e-05, 4.0935e-05, 4.3241e-05, 4.5563e-05, 4.7966e-05, 5.0369e-05, 
    5.2871e-05, 5.544e-05, 5.7896e-05, 6.025e-05, 6.2476e-05, 6.471e-05, 
    6.6568e-05, 6.8478e-05, 7.0319e-05, 7.1849e-05, 7.3166e-05, 7.4046e-05, 
    7.4634e-05, 7.5117e-05, 7.5459e-05, 7.5498e-05, 7.5177e-05, 7.4332e-05, 
    7.3068e-05, 7.1432e-05, 6.9399e-05, 6.6934e-05, 6.4046e-05, 6.1046e-05, 
    5.794e-05, 5.4791e-05, 5.1708e-05, 4.8809e-05, 4.6401e-05, 4.4275e-05, 
    4.2372e-05, 4.0584e-05, 3.9175e-05, 3.771e-05, 3.6328e-05, 3.4963e-05, 
    3.3446e-05, 3.1973e-05, 3.0539e-05, 2.9382e-05, 2.8484e-05, 2.7906e-05, 
    2.7827e-05, 2.8323e-05, 2.8726e-05, 2.981e-05, 3.0711e-05, 3.187e-05, 
    3.2948e-05, 3.4222e-05, 3.5677e-05, 3.7308e-05, 3.8744e-05, 4.0409e-05, 
    4.1909e-05, 4.3143e-05, 4.4384e-05, 4.5536e-05, 4.6621e-05, 4.77e-05, 
    4.8669e-05, 4.9465e-05, 5.0114e-05, 5.0206e-05, 4.9973e-05, 4.9519e-05, 
    4.8758e-05, 4.7369e-05, 4.5781e-05, 4.3931e-05, 4.176e-05, 3.9519e-05, 
    3.7024e-05, 3.4415e-05, 3.1865e-05, 2.9471e-05, 2.7163e-05, 2.4823e-05, 
    2.2656e-05, 2.0691e-05, 1.9341e-05, 1.8314e-05, 1.7684e-05, 1.726e-05, 
    1.6882e-05, 1.6427e-05, 1.5735e-05, 1.5027e-05, 1.4413e-05, 1.3977e-05, 
    1.4057e-05, 1.455e-05, 1.5484e-05, 1.7045e-05, 1.8672e-05, 2.0646e-05, 
    2.2856e-05, 2.492e-05, 2.6853e-05, 2.8627e-05, 3.0322e-05, 3.1867e-05, 
    3.3133e-05, 3.4201e-05, 3.5477e-05, 3.6458e-05, 3.7565e-05, 3.8252e-05, 
    3.9184e-05, 3.9826e-05, 4.0569e-05, 4.1512e-05, 4.2765e-05, 4.3898e-05, 
    4.5507e-05, 4.7185e-05, 4.8562e-05, 4.9817e-05, 5.0937e-05, 5.2065e-05, 
    5.3169e-05, 5.4303e-05, 5.5359e-05, 5.618e-05, 5.6841e-05, 5.752e-05, 
    5.8212e-05, 5.8794e-05, 5.9139e-05, 5.9482e-05, 5.9646e-05, 5.9486e-05, 
    5.93e-05, 5.8882e-05, 5.8108e-05, 5.7146e-05, 5.6007e-05, 5.442e-05, 
    5.2329e-05, 4.9936e-05, 4.7154e-05, 4.4315e-05, 4.1257e-05, 3.8327e-05, 
    3.5403e-05, 3.3001e-05, 3.0843e-05, 2.8594e-05, 2.6576e-05, 2.4865e-05, 
    2.3265e-05, 2.1984e-05, 2.1088e-05, 2.0783e-05, 2.1055e-05, 2.1558e-05, 
    2.2514e-05, 2.3778e-05, 2.5432e-05, 2.7237e-05, 2.9286e-05, 3.1491e-05, 
    3.3918e-05, 3.6383e-05, 3.8817e-05, 4.1203e-05, 4.3439e-05, 4.5358e-05, 
    4.6894e-05, 4.8074e-05, 4.8782e-05, 4.9008e-05, 4.8523e-05, 4.7788e-05, 
    4.6807e-05, 4.586e-05, 4.4937e-05, 4.3734e-05, 4.2373e-05, 4.0846e-05, 
    3.9311e-05, 3.7618e-05, 3.6067e-05, 3.4611e-05, 3.3171e-05, 3.1587e-05, 
    3.0247e-05, 2.9151e-05, 2.814e-05, 2.7215e-05, 2.6637e-05, 2.6228e-05, 
    2.615e-05, 2.6503e-05, 2.6978e-05, 2.7559e-05, 2.8333e-05, 2.951e-05, 
    3.0713e-05, 3.1827e-05, 3.2935e-05, 3.4092e-05, 3.5006e-05, 3.5819e-05, 
    3.6584e-05, 3.6841e-05, 3.7289e-05, 3.7626e-05, 3.7794e-05, 3.7778e-05, 
    3.7711e-05, 3.7265e-05, 3.6738e-05, 3.6048e-05, 3.539e-05, 3.4694e-05, 
    3.3897e-05, 3.3223e-05, 3.2439e-05, 3.1689e-05, 3.0922e-05, 3.0147e-05, 
    2.9361e-05, 2.8822e-05, 2.8413e-05, 2.8119e-05, 2.8079e-05, 2.8353e-05, 
    2.8836e-05, 2.9514e-05, 3.0471e-05, 3.1442e-05, 3.2403e-05, 3.3188e-05, 
    3.3811e-05, 3.4312e-05, 3.4862e-05, 3.5467e-05, 3.606e-05, 3.6572e-05, 
    3.7041e-05, 3.7357e-05, 3.7513e-05, 3.7625e-05, 3.7664e-05, 3.782e-05, 
    3.7762e-05, 3.7756e-05, 3.7566e-05, 3.7379e-05, 3.7279e-05, 3.7133e-05, 
    3.6899e-05, 3.6809e-05, 3.6819e-05, 3.6788e-05, 3.685e-05, 3.6954e-05, 
    3.7444e-05, 3.7854e-05, 3.8394e-05, 3.9122e-05, 4.0262e-05, 4.119e-05, 
    4.1999e-05, 4.2796e-05, 4.3309e-05, 4.4159e-05, 4.5191e-05, 4.6494e-05, 
    4.7814e-05, 4.9348e-05, 5.0387e-05, 5.1276e-05, 5.1775e-05, 5.2069e-05, 
    5.2021e-05, 5.1657e-05, 5.1167e-05, 5.0448e-05, 4.9571e-05, 4.8714e-05, 
    4.785e-05, 4.681e-05, 4.5809e-05, 4.4596e-05, 4.3378e-05, 4.2369e-05, 
    4.1466e-05, 4.0646e-05, 3.9931e-05, 3.9383e-05, 3.9139e-05, 3.8988e-05, 
    3.9394e-05, 4.0128e-05, 4.1171e-05, 4.2384e-05, 4.3941e-05, 4.5713e-05, 
    4.7551e-05, 4.9359e-05, 5.0995e-05, 5.2558e-05, 5.4007e-05, 5.5143e-05, 
    5.6098e-05, 5.6588e-05, 5.6799e-05, 5.6512e-05, 5.5772e-05, 5.4857e-05, 
    5.3447e-05, 5.1747e-05, 4.9855e-05, 4.7687e-05, 4.5367e-05, 4.2866e-05, 
    4.0194e-05, 3.767e-05, 3.4915e-05, 3.2071e-05, 2.9396e-05, 2.6877e-05, 
    2.4356e-05, 2.1739e-05, 1.8995e-05, 1.6021e-05, 1.341e-05, 1.1127e-05, 
    9.388e-06, 8.259e-06, 8.03e-06, 8.122e-06, 8.786e-06, 9.959e-06, 
    1.1279e-05, 1.3137e-05, 1.5312e-05, 1.7916e-05, 2.0847e-05, 2.391e-05, 
    2.6989e-05, 3.012e-05, 3.3046e-05, 3.5735e-05, 3.8138e-05, 4.0394e-05, 
    4.261e-05, 4.4548e-05, 4.6053e-05, 4.7315e-05, 4.813e-05, 4.8504e-05, 
    4.8191e-05, 4.7262e-05, 4.5855e-05, 4.3914e-05, 4.1677e-05, 3.9146e-05, 
    3.6508e-05, 3.3766e-05, 3.1212e-05, 2.8705e-05,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 0.002548, 0.0025362, 0.0025243, 
    0.0025124, 0.0025006, 0.0024887, 0.0024771, 0.0024656, 0.0024541, 
    0.0024431, 0.002432, 0.0024207, 0.0024094, 0.0023982, 0.002387, 
    0.0023757, 0.0023646, 0.0023533, 0.0023421, 0.0023309, 0.0023201, 
    0.0023093, 0.0022988, 0.0022881, 0.0022776, 0.0022668, 0.0022561, 
    0.0022454, 0.0022348, 0.0022246, 0.0022149, 0.002205, 0.0021955, 
    0.0021864, 0.0021776, 0.0021688, 0.0021598, 0.0021507, 0.0021414, 
    0.0021324, 0.0021231, 0.0021137, 0.0021044, 0.0020951, 0.002085, 
    0.0020751, 0.0020652, 0.0020548, 0.0020446, 0.002034, 0.0020235, 
    0.0020125, 0.0020016, 0.00199, 0.0019786, 0.0019668, 0.0019546, 
    0.0019426, 0.0019299, 0.0019176, 0.0019048, 0.001892, 0.0018789, 
    0.0018655, 0.001852, 0.0018387, 0.0018254, 0.0018125, 0.0017996, 
    0.0017869, 0.0017745, 0.0017626, 0.001751, 0.0017395, 0.0017287, 
    0.0017185, 0.0017082, 0.0016986, 0.0016895, 0.0016808, 0.0016722, 
    0.0016641, 0.0016563, 0.001649, 0.0016415, 0.0016347, 0.0016279, 
    0.0016212, 0.0016142, 0.0016077, 0.001601, 0.0015947, 0.0015879, 
    0.0015813, 0.0015746, 0.0015681, 0.0015617, 0.001555, 0.001548, 
    0.0015408, 0.0015341, 0.0015269, 0.0015196, 0.0015123, 0.001505, 
    0.0014972, 0.0014901, 0.0014826, 0.0014751, 0.0014678, 0.0014603, 
    0.0014528, 0.0014452, 0.0014376, 0.0014302, 0.0014228, 0.0014151, 
    0.0014076, 0.0014002, 0.0013924, 0.0013846, 0.0013768, 0.0013694, 
    0.0013616, 0.0013537, 0.001346, 0.001338, 0.0013301, 0.0013222, 
    0.0013142, 0.0013063, 0.0012981, 0.0012901, 0.0012818, 0.0012735, 
    0.0012651, 0.0012568, 0.0012483, 0.0012401, 0.001232, 0.0012239, 
    0.0012156, 0.0012076, 0.0011995, 0.0011914, 0.0011831, 0.0011749, 
    0.0011669, 0.0011589, 0.0011509, 0.0011433, 0.0011356, 0.0011279, 
    0.0011205, 0.001113, 0.0011058, 0.0010986, 0.0010916, 0.0010847, 
    0.0010777, 0.0010706, 0.0010642, 0.0010573, 0.0010509, 0.0010447, 
    0.0010385, 0.0010323, 0.0010265, 0.0010209, 0.0010153, 0.0010099, 
    0.0010047, 0.00099967, 0.00099492, 0.00099023, 0.00098577, 0.00098165, 
    0.00097747, 0.00097346, 0.00096921, 0.00096496, 0.00096071, 0.0009564, 
    0.00095231, 0.00094779, 0.00094328, 0.0009388, 0.00093422, 0.00092929, 
    0.00092443, 0.00091934, 0.00091422, 0.00090894, 0.00090347, 0.00089762, 
    0.00089163, 0.00088509, 0.00087858, 0.0008716, 0.00086489, 0.00085803, 
    0.00085102, 0.00084392, 0.00083687, 0.00082974, 0.00082257, 0.0008152, 
    0.00080763, 0.00080024, 0.00079265, 0.00078513, 0.00077787, 0.00077059, 
    0.0007635, 0.0007567, 0.00074981, 0.00074344, 0.00073712, 0.0007311, 
    0.00072531, 0.00071978, 0.00071419, 0.00070906, 0.00070418, 0.0006995, 
    0.00069486, 0.00069081, 0.00068675, 0.0006829, 0.00067922, 0.00067555, 
    0.0006719, 0.00066822, 0.00066453, 0.00066098, 0.00065716, 0.00065331, 
    0.00064953, 0.00064572, 0.00064166, 0.00063712, 0.00063229, 0.00062743, 
    0.00062256, 0.00061757, 0.00061229, 0.00060709, 0.00060163, 0.00059629, 
    0.0005908, 0.00058549, 0.00058026, 0.00057507, 0.00056996, 0.00056498, 
    0.00056028, 0.00055557, 0.00055082, 0.00054615, 0.00054163, 0.00053717, 
    0.00053289, 0.00052852, 0.00052446, 0.00052065, 0.00051692, 0.00051349, 
    0.00051022, 0.00050712, 0.00050424, 0.00050153, 0.00049888, 0.00049618, 
    0.00049333, 0.00049071, 0.00048821, 0.00048562, 0.00048291, 0.00048012, 
    0.00047719, 0.00047399, 0.00047086, 0.00046773, 0.00046458, 0.00046141, 
    0.00045783, 0.00045394, 0.0004503, 0.00044647, 0.00044264, 0.00043889, 
    0.00043517, 0.00043144, 0.00042792, 0.0004245, 0.00042126, 0.00041787, 
    0.00041468, 0.00041159, 0.00040852, 0.00040545, 0.00040245, 0.00039948, 
    0.00039674, 0.00039429, 0.00039192, 0.0003894, 0.00038736, 0.00038523, 
    0.00038307, 0.00038098, 0.00037883, 0.00037665, 0.00037449, 0.00037215, 
    0.00037003, 0.00036803, 0.00036616, 0.00036463, 0.00036301, 0.00036162, 
    0.00036029, 0.00035902, 0.0003578, 0.00035662, 0.00035532, 0.00035394, 
    0.00035249, 0.000351, 0.0003495, 0.00034789, 0.00034628, 0.00034491, 
    0.00034355, 0.00034196, 0.00034038, 0.00033873, 0.00033711, 0.00033538, 
    0.00033371, 0.0003317, 0.00032935, 0.00032688, 0.00032438, 0.00032182, 
    0.00031905, 0.00031606, 0.00031303, 0.00030986, 0.0003064, 0.00030289, 
    0.00029923, 0.00029527, 0.00029133, 0.0002875, 0.00028364, 0.00027992, 
    0.00027622, 0.00027265, 0.00026911, 0.0002658, 0.00026225, 0.0002588, 
    0.00025548, 0.00025222, 0.00024912, 0.00024634, 0.0002436, 0.00024123, 
    0.00023919, 0.00023742, 0.00023573, 0.00023435, 0.00023305, 0.00023188, 
    0.00023072, 0.00022962, 0.00022856, 0.00022752, 0.00022666, 0.00022579, 
    0.00022488, 0.00022413, 0.00022336, 0.00022288, 0.00022234, 0.00022185, 
    0.00022116, 0.00022036, 0.00021949, 0.00021853, 0.00021723, 0.00021562, 
    0.00021411, 0.00021263, 0.00021081, 0.00020896, 0.00020718, 0.00020532, 
    0.00020352, 0.00020196, 0.00020014, 0.00019844, 0.00019676, 0.00019512, 
    0.00019364, 0.00019217, 0.00019085, 0.00018973, 0.0001887, 0.00018772, 
    0.00018687, 0.0001862, 0.00018534, 0.00018464, 0.0001839, 0.00018335, 
    0.00018283, 0.00018235, 0.0001817, 0.000181, 0.00018065, 0.00017997, 
    0.00017915, 0.00017841, 0.00017771, 0.00017679, 0.00017577, 0.00017452, 
    0.0001729, 0.00017133, 0.00016966, 0.00016777, 0.00016597, 0.00016427, 
    0.00016245, 0.00016059, 0.00015877, 0.00015707, 0.00015532, 0.00015359, 
    0.0001518, 0.00015008, 0.00014845, 0.00014673, 0.00014521, 0.00014383, 
    0.00014263, 0.00014139, 0.00014022, 0.0001392, 0.00013844, 0.00013763, 
    0.00013687, 0.00013622, 0.00013565, 0.00013516, 0.00013475, 0.00013424, 
    0.00013373, 0.00013325, 0.00013288, 0.0001322, 0.00013155, 0.00013088, 
    0.00013007, 0.00012929, 0.00012847, 0.0001275, 0.00012645, 0.00012513, 
    0.00012375, 0.00012233, 0.00012076, 0.00011932, 0.0001178, 0.00011578, 
    0.00011418, 0.00011263, 0.00011121, 0.00010966, 0.0001082, 0.00010696, 
    0.0001056, 0.00010405, 0.00010262, 0.00010139, 0.00010028, 9.9289e-05, 
    9.8352e-05, 9.7269e-05, 9.6322e-05, 9.5355e-05, 9.4581e-05, 9.3888e-05, 
    9.3395e-05, 9.2822e-05, 9.2375e-05, 9.215e-05, 9.2274e-05, 9.2429e-05, 
    9.2745e-05, 9.3209e-05, 9.4e-05, 9.4923e-05, 9.5877e-05, 9.6805e-05, 
    9.789e-05, 9.9109e-05, 0.00010036, 0.00010156, 0.00010263, 0.00010375, 
    0.00010442, 0.00010514, 0.00010561, 0.00010587, 0.00010605, 0.00010631, 
    0.00010637, 0.00010625, 0.00010592, 0.00010546, 0.00010479, 0.00010427, 
    0.00010375, 0.00010294, 0.00010221, 0.00010131, 0.00010035, 9.9014e-05, 
    9.7613e-05, 9.5878e-05, 9.4195e-05, 9.2275e-05, 9.0662e-05, 8.895e-05, 
    8.6734e-05, 8.4683e-05, 8.26e-05, 8.0543e-05, 7.855e-05, 7.6785e-05, 
    7.5073e-05, 7.3427e-05, 7.1873e-05, 7.0415e-05, 6.8886e-05, 6.7577e-05, 
    6.6443e-05, 6.5413e-05, 6.4427e-05, 6.3657e-05, 6.2924e-05, 6.2247e-05, 
    6.1582e-05, 6.1078e-05, 6.0515e-05, 5.9845e-05, 5.9185e-05, 5.8599e-05, 
    5.779e-05, 5.7125e-05, 5.6364e-05, 5.5719e-05, 5.5069e-05, 5.4394e-05, 
    5.3517e-05, 5.2559e-05, 5.1677e-05, 5.0936e-05, 5.0524e-05, 5.012e-05, 
    4.9927e-05, 4.9543e-05, 4.9397e-05, 4.9436e-05, 4.9263e-05, 4.9199e-05, 
    4.9321e-05, 4.9631e-05, 4.9917e-05, 5.0107e-05, 5.0077e-05, 5.0002e-05, 
    5.0148e-05, 5.0411e-05, 5.0464e-05, 5.0892e-05, 5.1089e-05, 5.1535e-05, 
    5.1743e-05, 5.222e-05, 5.2405e-05, 5.2622e-05, 5.2804e-05, 5.3277e-05, 
    5.3783e-05, 5.4235e-05, 5.4696e-05, 5.5105e-05, 5.5316e-05, 5.551e-05, 
    5.5772e-05, 5.5965e-05, 5.6215e-05, 5.6583e-05, 5.6922e-05, 5.6966e-05, 
    5.6919e-05, 5.6883e-05, 5.6578e-05, 5.6111e-05, 5.5599e-05, 5.4976e-05, 
    5.4225e-05, 5.3386e-05, 5.2707e-05, 5.2233e-05, 5.1704e-05, 5.1392e-05, 
    5.1276e-05, 5.1244e-05, 5.1634e-05, 5.2083e-05, 5.2729e-05, 5.3195e-05, 
    5.4194e-05, 5.5603e-05, 5.7075e-05, 5.8722e-05, 6.061e-05, 6.2878e-05, 
    6.5221e-05, 6.7812e-05, 7.0325e-05, 7.2923e-05, 7.5713e-05, 7.8212e-05, 
    8.0591e-05, 8.2984e-05, 8.4986e-05, 8.6869e-05, 8.8362e-05, 8.9439e-05, 
    9.0055e-05, 9.0312e-05, 9.0199e-05, 8.9608e-05, 8.8774e-05, 8.7384e-05, 
    8.5764e-05, 8.376e-05, 8.1353e-05, 7.858e-05, 7.5539e-05, 7.2238e-05, 
    6.8849e-05, 6.5368e-05, 6.178e-05, 5.8019e-05, 5.4237e-05, 5.0365e-05, 
    4.6464e-05, 4.2652e-05, 3.9075e-05, 3.5674e-05, 3.2772e-05, 3.0385e-05, 
    2.8111e-05, 2.6242e-05, 2.4846e-05, 2.3637e-05, 2.2767e-05, 2.244e-05, 
    2.2163e-05, 2.2242e-05, 2.2549e-05, 2.308e-05, 2.3761e-05, 2.4746e-05, 
    2.6e-05, 2.7325e-05, 2.9055e-05, 3.1064e-05, 3.3104e-05, 3.5222e-05, 
    3.6899e-05, 3.8647e-05, 4.0339e-05, 4.1715e-05, 4.3029e-05, 4.4071e-05, 
    4.5131e-05, 4.5894e-05, 4.6569e-05, 4.7012e-05, 4.7246e-05, 4.7269e-05, 
    4.7193e-05, 4.6902e-05, 4.6736e-05, 4.6118e-05, 4.5441e-05, 4.4553e-05, 
    4.3532e-05, 4.2481e-05, 4.1169e-05, 3.9896e-05, 3.8586e-05, 3.731e-05, 
    3.5973e-05, 3.4791e-05, 3.3834e-05, 3.2878e-05, 3.1954e-05, 3.1029e-05, 
    3.0196e-05, 2.935e-05, 2.8771e-05, 2.8273e-05, 2.7869e-05, 2.7455e-05, 
    2.7197e-05, 2.6952e-05, 2.6764e-05, 2.6718e-05, 2.6693e-05, 2.6903e-05, 
    2.7309e-05, 2.7876e-05, 2.8471e-05, 2.9398e-05, 3.0578e-05, 3.1815e-05, 
    3.336e-05, 3.4804e-05, 3.644e-05, 3.8328e-05, 4.0526e-05, 4.273e-05, 
    4.5081e-05, 4.7109e-05, 4.8886e-05, 5.0451e-05, 5.166e-05, 5.2413e-05, 
    5.2758e-05, 5.2847e-05, 5.2737e-05, 5.2246e-05, 5.1466e-05, 5.0629e-05, 
    4.9596e-05, 4.8561e-05, 4.7453e-05, 4.6371e-05, 4.5223e-05, 4.4252e-05, 
    4.3123e-05, 4.1988e-05, 4.1053e-05, 4.034e-05, 3.9921e-05, 3.9544e-05, 
    3.9698e-05, 3.9895e-05, 4.0319e-05, 4.0806e-05, 4.1462e-05, 4.228e-05, 
    4.3146e-05, 4.3931e-05, 4.4797e-05, 4.5575e-05, 4.6466e-05, 4.7333e-05, 
    4.8102e-05, 4.8801e-05, 4.9353e-05, 4.9964e-05, 5.057e-05, 5.1119e-05, 
    5.1545e-05, 5.1936e-05, 5.2105e-05, 5.2046e-05, 5.178e-05, 5.1311e-05, 
    5.077e-05, 5.0173e-05, 4.9453e-05, 4.8351e-05, 4.7072e-05, 4.5809e-05, 
    4.4298e-05, 4.2453e-05, 4.0055e-05, 3.7445e-05, 3.459e-05, 3.1961e-05, 
    2.9494e-05, 2.7145e-05, 2.4905e-05, 2.322e-05, 2.1831e-05, 2.0849e-05, 
    2.0119e-05, 1.9498e-05, 1.9124e-05, 1.8659e-05, 1.8586e-05, 1.8453e-05, 
    1.8694e-05, 1.9119e-05, 1.9632e-05, 2.0372e-05, 2.1282e-05, 2.2291e-05, 
    2.3645e-05, 2.4927e-05, 2.6117e-05, 2.7361e-05, 2.8138e-05, 2.8941e-05, 
    2.931e-05, 2.9892e-05, 3.0269e-05, 3.0473e-05, 3.0995e-05, 3.1212e-05, 
    3.1405e-05, 3.1492e-05, 3.138e-05, 3.1295e-05, 3.0839e-05, 3.0424e-05, 
    2.9853e-05, 2.9283e-05, 2.8562e-05, 2.7923e-05, 2.7319e-05, 2.7004e-05, 
    2.6725e-05, 2.647e-05, 2.6549e-05, 2.6697e-05, 2.6838e-05, 2.7158e-05, 
    2.7204e-05, 2.7112e-05, 2.7352e-05, 2.757e-05, 2.7867e-05, 2.8216e-05, 
    2.8964e-05, 2.9958e-05, 3.1267e-05, 3.2757e-05, 3.455e-05, 3.6442e-05, 
    3.8544e-05, 4.0935e-05, 4.3241e-05, 4.5563e-05, 4.7966e-05, 5.0369e-05, 
    5.2871e-05, 5.544e-05, 5.7896e-05, 6.025e-05, 6.2476e-05, 6.471e-05, 
    6.6568e-05, 6.8478e-05, 7.0319e-05, 7.1849e-05, 7.3166e-05, 7.4046e-05, 
    7.4634e-05, 7.5117e-05, 7.5459e-05, 7.5498e-05, 7.5177e-05, 7.4332e-05, 
    7.3068e-05, 7.1432e-05, 6.9399e-05, 6.6934e-05, 6.4046e-05, 6.1046e-05, 
    5.794e-05, 5.4791e-05, 5.1708e-05, 4.8809e-05, 4.6401e-05, 4.4275e-05, 
    4.2372e-05, 4.0584e-05, 3.9175e-05, 3.771e-05, 3.6328e-05, 3.4963e-05, 
    3.3446e-05, 3.1973e-05, 3.0539e-05, 2.9382e-05, 2.8484e-05, 2.7906e-05, 
    2.7827e-05, 2.8323e-05, 2.8726e-05, 2.981e-05, 3.0711e-05, 3.187e-05, 
    3.2948e-05, 3.4222e-05, 3.5677e-05, 3.7308e-05, 3.8744e-05, 4.0409e-05, 
    4.1909e-05, 4.3143e-05, 4.4384e-05, 4.5536e-05, 4.6621e-05, 4.77e-05, 
    4.8669e-05, 4.9465e-05, 5.0114e-05, 5.0206e-05, 4.9973e-05, 4.9519e-05, 
    4.8758e-05, 4.7369e-05, 4.5781e-05, 4.3931e-05, 4.176e-05, 3.9519e-05, 
    3.7024e-05, 3.4415e-05, 3.1865e-05, 2.9471e-05, 2.7163e-05, 2.4823e-05, 
    2.2656e-05, 2.0691e-05, 1.9341e-05, 1.8314e-05, 1.7684e-05, 1.726e-05, 
    1.6882e-05, 1.6427e-05, 1.5735e-05, 1.5027e-05, 1.4413e-05, 1.3977e-05, 
    1.4057e-05, 1.455e-05, 1.5484e-05, 1.7045e-05, 1.8672e-05, 2.0646e-05, 
    2.2856e-05, 2.492e-05, 2.6853e-05, 2.8627e-05, 3.0322e-05, 3.1867e-05, 
    3.3133e-05, 3.4201e-05, 3.5477e-05, 3.6458e-05, 3.7565e-05, 3.8252e-05, 
    3.9184e-05, 3.9826e-05, 4.0569e-05, 4.1512e-05, 4.2765e-05, 4.3898e-05, 
    4.5507e-05, 4.7185e-05, 4.8562e-05, 4.9817e-05, 5.0937e-05, 5.2065e-05, 
    5.3169e-05, 5.4303e-05, 5.5359e-05, 5.618e-05, 5.6841e-05, 5.752e-05, 
    5.8212e-05, 5.8794e-05, 5.9139e-05, 5.9482e-05, 5.9646e-05, 5.9486e-05, 
    5.93e-05, 5.8882e-05, 5.8108e-05, 5.7146e-05, 5.6007e-05, 5.442e-05, 
    5.2329e-05, 4.9936e-05, 4.7154e-05, 4.4315e-05, 4.1257e-05, 3.8327e-05, 
    3.5403e-05, 3.3001e-05, 3.0843e-05, 2.8594e-05, 2.6576e-05, 2.4865e-05, 
    2.3265e-05, 2.1984e-05, 2.1088e-05, 2.0783e-05, 2.1055e-05, 2.1558e-05, 
    2.2514e-05, 2.3778e-05, 2.5432e-05, 2.7237e-05, 2.9286e-05, 3.1491e-05, 
    3.3918e-05, 3.6383e-05, 3.8817e-05, 4.1203e-05, 4.3439e-05, 4.5358e-05, 
    4.6894e-05, 4.8074e-05, 4.8782e-05, 4.9008e-05, 4.8523e-05, 4.7788e-05, 
    4.6807e-05, 4.586e-05, 4.4937e-05, 4.3734e-05, 4.2373e-05, 4.0846e-05, 
    3.9311e-05, 3.7618e-05, 3.6067e-05, 3.4611e-05, 3.3171e-05, 3.1587e-05, 
    3.0247e-05, 2.9151e-05, 2.814e-05, 2.7215e-05, 2.6637e-05, 2.6228e-05, 
    2.615e-05, 2.6503e-05, 2.6978e-05, 2.7559e-05, 2.8333e-05, 2.951e-05, 
    3.0713e-05, 3.1827e-05, 3.2935e-05, 3.4092e-05, 3.5006e-05, 3.5819e-05, 
    3.6584e-05, 3.6841e-05, 3.7289e-05, 3.7626e-05, 3.7794e-05, 3.7778e-05, 
    3.7711e-05, 3.7265e-05, 3.6738e-05, 3.6048e-05, 3.539e-05, 3.4694e-05, 
    3.3897e-05, 3.3223e-05, 3.2439e-05, 3.1689e-05, 3.0922e-05, 3.0147e-05, 
    2.9361e-05, 2.8822e-05, 2.8413e-05, 2.8119e-05, 2.8079e-05, 2.8353e-05, 
    2.8836e-05, 2.9514e-05, 3.0471e-05, 3.1442e-05, 3.2403e-05, 3.3188e-05, 
    3.3811e-05, 3.4312e-05, 3.4862e-05, 3.5467e-05, 3.606e-05, 3.6572e-05, 
    3.7041e-05, 3.7357e-05, 3.7513e-05, 3.7625e-05, 3.7664e-05, 3.782e-05, 
    3.7762e-05, 3.7756e-05, 3.7566e-05, 3.7379e-05, 3.7279e-05, 3.7133e-05, 
    3.6899e-05, 3.6809e-05, 3.6819e-05, 3.6788e-05, 3.685e-05, 3.6954e-05, 
    3.7444e-05, 3.7854e-05, 3.8394e-05, 3.9122e-05, 4.0262e-05, 4.119e-05, 
    4.1999e-05, 4.2796e-05, 4.3309e-05, 4.4159e-05, 4.5191e-05, 4.6494e-05, 
    4.7814e-05, 4.9348e-05, 5.0387e-05, 5.1276e-05, 5.1775e-05, 5.2069e-05, 
    5.2021e-05, 5.1657e-05, 5.1167e-05, 5.0448e-05, 4.9571e-05, 4.8714e-05, 
    4.785e-05, 4.681e-05, 4.5809e-05, 4.4596e-05, 4.3378e-05, 4.2369e-05, 
    4.1466e-05, 4.0646e-05, 3.9931e-05, 3.9383e-05, 3.9139e-05, 3.8988e-05, 
    3.9394e-05, 4.0128e-05, 4.1171e-05, 4.2384e-05, 4.3941e-05, 4.5713e-05, 
    4.7551e-05, 4.9359e-05, 5.0995e-05, 5.2558e-05, 5.4007e-05, 5.5143e-05, 
    5.6098e-05, 5.6588e-05, 5.6799e-05, 5.6512e-05, 5.5772e-05, 5.4857e-05, 
    5.3447e-05, 5.1747e-05, 4.9855e-05, 4.7687e-05, 4.5367e-05, 4.2866e-05, 
    4.0194e-05, 3.767e-05, 3.4915e-05, 3.2071e-05, 2.9396e-05, 2.6877e-05, 
    2.4356e-05, 2.1739e-05, 1.8995e-05, 1.6021e-05, 1.341e-05, 1.1127e-05, 
    9.388e-06, 8.259e-06, 8.03e-06, 8.122e-06, 8.786e-06, 9.959e-06, 
    1.1279e-05, 1.3137e-05, 1.5312e-05, 1.7916e-05, 2.0847e-05, 2.391e-05, 
    2.6989e-05, 3.012e-05, 3.3046e-05, 3.5735e-05, 3.8138e-05, 4.0394e-05, 
    4.261e-05, 4.4548e-05, 4.6053e-05, 4.7315e-05, 4.813e-05, 4.8504e-05, 
    4.8191e-05, 4.7262e-05, 4.5855e-05, 4.3914e-05, 4.1677e-05, 3.9146e-05, 
    3.6508e-05, 3.3766e-05, 3.1212e-05, 2.8705e-05 ;

 bangle =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 0.0021696, 0.0021573, 0.0021454, 
    0.0021335, 0.0021214, 0.0021092, 0.0020971, 0.0020854, 0.0020741, 
    0.002063, 0.0020521, 0.0020412, 0.0020307, 0.0020203, 0.0020099, 
    0.0019995, 0.0019901, 0.0019804, 0.0019709, 0.0019621, 0.0019529, 
    0.0019446, 0.0019365, 0.0019288, 0.0019218, 0.0019149, 0.0019084, 
    0.0019028, 0.0018967, 0.0018919, 0.0018871, 0.0018827, 0.0018789, 
    0.0018763, 0.0018732, 0.0018691, 0.0018637, 0.001858, 0.0018513, 
    0.0018435, 0.0018348, 0.0018258, 0.001816, 0.0018054, 0.0017945, 
    0.0017833, 0.0017717, 0.0017598, 0.001748, 0.0017363, 0.0017246, 
    0.0017131, 0.0017016, 0.0016906, 0.0016793, 0.0016683, 0.0016574, 
    0.0016469, 0.0016364, 0.0016259, 0.0016155, 0.0016053, 0.0015953, 
    0.0015853, 0.0015754, 0.0015655, 0.0015556, 0.0015458, 0.0015363, 
    0.0015269, 0.0015173, 0.0015078, 0.0014986, 0.0014894, 0.0014802, 
    0.0014712, 0.0014621, 0.0014529, 0.0014439, 0.0014348, 0.0014258, 
    0.0014169, 0.0014082, 0.0013996, 0.0013911, 0.0013828, 0.0013744, 
    0.0013665, 0.0013586, 0.0013508, 0.0013434, 0.0013362, 0.0013292, 
    0.001322, 0.0013152, 0.0013085, 0.0013019, 0.0012956, 0.0012893, 
    0.0012832, 0.001277, 0.001271, 0.0012652, 0.0012595, 0.0012539, 
    0.0012483, 0.0012426, 0.0012369, 0.0012307, 0.0012242, 0.0012176, 
    0.0012111, 0.0012042, 0.0011971, 0.00119, 0.001183, 0.0011759, 0.0011684, 
    0.0011609, 0.0011533, 0.0011452, 0.0011372, 0.0011292, 0.0011211, 
    0.001113, 0.0011047, 0.0010966, 0.0010886, 0.0010806, 0.001073, 
    0.0010656, 0.0010581, 0.001051, 0.001044, 0.0010371, 0.0010305, 
    0.0010242, 0.0010178, 0.0010116, 0.0010057, 0.00099995, 0.0009944, 
    0.00098904, 0.00098375, 0.00097859, 0.00097346, 0.00096835, 0.0009633, 
    0.0009582, 0.00095317, 0.00094811, 0.00094303, 0.00093786, 0.00093253, 
    0.00092711, 0.0009216, 0.00091593, 0.00091006, 0.00090409, 0.00089794, 
    0.0008916, 0.00088503, 0.00087825, 0.00087138, 0.00086437, 0.00085731, 
    0.00085019, 0.00084312, 0.00083595, 0.00082885, 0.00082148, 0.00081415, 
    0.00080699, 0.00079992, 0.00079284, 0.00078585, 0.00077893, 0.00077234, 
    0.000766, 0.00075973, 0.00075371, 0.00074774, 0.00074182, 0.00073604, 
    0.00073031, 0.00072466, 0.00071909, 0.00071351, 0.00070805, 0.00070259, 
    0.00069721, 0.00069202, 0.00068692, 0.00068183, 0.00067677, 0.00067184, 
    0.00066691, 0.00066199, 0.00065709, 0.00065221, 0.00064737, 0.0006426, 
    0.00063792, 0.00063329, 0.0006287, 0.00062413, 0.00061965, 0.00061522, 
    0.00061077, 0.00060635, 0.00060205, 0.00059786, 0.0005938, 0.00058971, 
    0.00058566, 0.00058168, 0.00057777, 0.00057394, 0.00057019, 0.00056655, 
    0.00056301, 0.00055949, 0.00055601, 0.00055251, 0.000549, 0.0005454, 
    0.0005418, 0.00053824, 0.00053468, 0.00053111, 0.00052756, 0.00052397, 
    0.00052042, 0.00051685, 0.00051326, 0.00050969, 0.0005061, 0.00050249, 
    0.0004989, 0.00049533, 0.00049175, 0.00048818, 0.00048464, 0.00048113, 
    0.00047758, 0.00047398, 0.00047036, 0.00046677, 0.00046319, 0.00045964, 
    0.00045615, 0.00045263, 0.00044912, 0.00044559, 0.00044206, 0.00043854, 
    0.0004351, 0.00043163, 0.00042814, 0.00042467, 0.00042115, 0.00041764, 
    0.00041418, 0.00041069, 0.00040723, 0.00040376, 0.00040036, 0.00039703, 
    0.00039372, 0.00039048, 0.00038732, 0.00038424, 0.0003812, 0.00037819, 
    0.00037517, 0.00037217, 0.00036926, 0.00036638, 0.0003635, 0.00036068, 
    0.0003579, 0.00035516, 0.00035247, 0.00034983, 0.00034721, 0.0003446, 
    0.00034198, 0.00033937, 0.00033675, 0.00033412, 0.00033152, 0.00032893, 
    0.00032637, 0.00032382, 0.00032128, 0.00031877, 0.00031628, 0.00031382, 
    0.00031139, 0.00030899, 0.00030661, 0.00030425, 0.00030191, 0.00029957, 
    0.00029722, 0.00029491, 0.0002926, 0.00029028, 0.00028794, 0.00028561, 
    0.00028326, 0.00028097, 0.00027875, 0.00027654, 0.00027434, 0.00027214, 
    0.00026995, 0.00026779, 0.0002656, 0.00026343, 0.00026132, 0.0002592, 
    0.00025711, 0.00025508, 0.00025301, 0.00025092, 0.0002488, 0.00024663, 
    0.00024448, 0.00024231, 0.00024014, 0.00023799, 0.00023591, 0.00023387, 
    0.00023183, 0.00022982, 0.00022778, 0.00022574, 0.00022371, 0.00022167, 
    0.00021966, 0.0002177, 0.00021578, 0.0002139, 0.00021208, 0.00021031, 
    0.00020856, 0.00020687, 0.00020522, 0.0002036, 0.00020202, 0.00020048, 
    0.00019896, 0.00019745, 0.00019594, 0.00019443, 0.00019292, 0.00019142, 
    0.00018992, 0.00018841, 0.00018692, 0.00018544, 0.00018399, 0.00018255, 
    0.00018111, 0.00017966, 0.00017822, 0.00017677, 0.00017532, 0.00017389, 
    0.00017244, 0.00017102, 0.00016964, 0.00016828, 0.00016693, 0.0001656, 
    0.00016428, 0.00016299, 0.00016171, 0.00016044, 0.0001592, 0.00015798, 
    0.00015677, 0.00015559, 0.00015442, 0.00015325, 0.00015208, 0.00015091, 
    0.00014973, 0.00014856, 0.0001474, 0.00014624, 0.00014508, 0.00014393, 
    0.00014279, 0.00014164, 0.0001405, 0.00013936, 0.00013821, 0.00013711, 
    0.00013602, 0.00013494, 0.00013388, 0.00013284, 0.00013179, 0.00013075, 
    0.00012973, 0.0001287, 0.00012765, 0.00012661, 0.00012556, 0.00012454, 
    0.00012352, 0.00012252, 0.00012153, 0.00012053, 0.00011954, 0.00011853, 
    0.00011753, 0.00011652, 0.00011551, 0.00011449, 0.00011347, 0.00011246, 
    0.00011145, 0.00011045, 0.00010945, 0.00010844, 0.00010744, 0.00010644, 
    0.00010545, 0.00010446, 0.00010347, 0.0001025, 0.00010154, 0.00010058, 
    9.9631e-05, 9.8686e-05, 9.7742e-05, 9.6814e-05, 9.5899e-05, 9.501e-05, 
    9.4148e-05, 9.3298e-05, 9.2462e-05, 9.1631e-05, 9.0856e-05, 9.0102e-05, 
    8.933e-05, 8.8552e-05, 8.7777e-05, 8.7006e-05, 8.6229e-05, 8.5462e-05, 
    8.4724e-05, 8.3997e-05, 8.3237e-05, 8.2457e-05, 8.1649e-05, 8.0825e-05, 
    8.001e-05, 7.9192e-05, 7.8386e-05, 7.7583e-05, 7.6781e-05, 7.5974e-05, 
    7.5176e-05, 7.4386e-05, 7.3609e-05, 7.2852e-05, 7.2123e-05, 7.1421e-05, 
    7.0745e-05, 7.0108e-05, 6.9496e-05, 6.8908e-05, 6.8338e-05, 6.7786e-05, 
    6.7264e-05, 6.6766e-05, 6.6283e-05, 6.5818e-05, 6.536e-05, 6.4899e-05, 
    6.4426e-05, 6.3955e-05, 6.3464e-05, 6.2965e-05, 6.2465e-05, 6.1967e-05, 
    6.1457e-05, 6.0941e-05, 6.0417e-05, 5.9882e-05, 5.9339e-05, 5.8783e-05, 
    5.8223e-05, 5.7679e-05, 5.7124e-05, 5.6564e-05, 5.6016e-05, 5.5503e-05, 
    5.4996e-05, 5.4532e-05, 5.4056e-05, 5.3599e-05, 5.3114e-05, 5.2668e-05, 
    5.2295e-05, 5.191e-05, 5.1541e-05, 5.118e-05, 5.0801e-05, 5.0415e-05, 
    5.0034e-05, 4.966e-05, 4.9297e-05, 4.8943e-05, 4.8587e-05, 4.8225e-05, 
    4.7859e-05, 4.7498e-05, 4.7138e-05, 4.6792e-05, 4.6447e-05, 4.6107e-05, 
    4.5761e-05, 4.5422e-05, 4.5084e-05, 4.4741e-05, 4.4395e-05, 4.4057e-05, 
    4.371e-05, 4.3365e-05, 4.3014e-05, 4.2656e-05, 4.2294e-05, 4.1951e-05, 
    4.1609e-05, 4.1261e-05, 4.0908e-05, 4.0552e-05, 4.0199e-05, 3.985e-05, 
    3.951e-05, 3.9165e-05, 3.8816e-05, 3.8469e-05, 3.8131e-05, 3.7808e-05, 
    3.7498e-05, 3.7207e-05, 3.6917e-05, 3.6625e-05, 3.6328e-05, 3.6027e-05, 
    3.5725e-05, 3.5422e-05, 3.5118e-05, 3.4811e-05, 3.4513e-05, 3.4212e-05, 
    3.3914e-05, 3.3615e-05, 3.331e-05, 3.3018e-05, 3.2761e-05, 3.254e-05, 
    3.2336e-05, 3.2143e-05, 3.1954e-05, 3.1765e-05, 3.1569e-05, 3.1367e-05, 
    3.116e-05, 3.0945e-05, 3.0717e-05, 3.047e-05, 3.0205e-05, 2.9928e-05, 
    2.9638e-05, 2.9347e-05, 2.9063e-05, 2.8788e-05, 2.8522e-05, 2.8262e-05, 
    2.8015e-05, 2.7783e-05, 2.7554e-05, 2.7329e-05, 2.7109e-05, 2.6894e-05, 
    2.668e-05, 2.6473e-05, 2.6284e-05, 2.6093e-05, 2.5896e-05, 2.5689e-05, 
    2.5518e-05, 2.5369e-05, 2.5224e-05, 2.5096e-05, 2.5005e-05, 2.4945e-05, 
    2.489e-05, 2.4849e-05, 2.4793e-05, 2.4748e-05, 2.4729e-05, 2.4658e-05, 
    2.4577e-05, 2.4489e-05, 2.4339e-05, 2.4139e-05, 2.3847e-05, 2.3458e-05, 
    2.2975e-05, 2.2419e-05, 2.1803e-05, 2.1151e-05, 2.0492e-05, 1.9852e-05, 
    1.9248e-05, 1.8704e-05, 1.8245e-05, 1.7891e-05, 1.7642e-05, 1.7519e-05, 
    1.7535e-05, 1.7648e-05, 1.7887e-05, 1.8239e-05, 1.8661e-05, 1.912e-05, 
    1.9594e-05, 2.0014e-05, 2.0309e-05, 2.0484e-05, 2.0523e-05, 2.0516e-05, 
    2.045e-05, 2.0319e-05, 2.0143e-05, 1.9918e-05, 1.9672e-05, 1.9428e-05, 
    1.9191e-05, 1.8978e-05, 1.8798e-05, 1.8641e-05, 1.8529e-05, 1.8457e-05, 
    1.8411e-05, 1.8412e-05, 1.8448e-05, 1.8508e-05, 1.8571e-05, 1.8608e-05, 
    1.8602e-05, 1.8575e-05, 1.8491e-05, 1.8357e-05, 1.818e-05, 1.7966e-05, 
    1.7712e-05, 1.7408e-05, 1.706e-05, 1.6678e-05, 1.6279e-05, 1.5889e-05, 
    1.5526e-05, 1.5194e-05, 1.4893e-05, 1.4627e-05, 1.4394e-05, 1.4201e-05, 
    1.4057e-05, 1.396e-05, 1.3916e-05, 1.3872e-05, 1.3848e-05, 1.3828e-05, 
    1.381e-05, 1.3786e-05, 1.3756e-05, 1.3734e-05, 1.3715e-05, 1.3697e-05, 
    1.3661e-05, 1.3607e-05, 1.3547e-05, 1.3491e-05, 1.3441e-05, 1.3389e-05, 
    1.3343e-05, 1.33e-05, 1.3257e-05, 1.3225e-05, 1.3192e-05, 1.3161e-05, 
    1.3136e-05, 1.3096e-05, 1.305e-05, 1.2999e-05, 1.2938e-05, 1.2867e-05, 
    1.2771e-05, 1.267e-05, 1.2584e-05, 1.2524e-05, 1.248e-05, 1.2439e-05, 
    1.2376e-05, 1.2271e-05, 1.2134e-05, 1.1979e-05, 1.1808e-05, 1.1633e-05, 
    1.1461e-05, 1.1306e-05, 1.1165e-05, 1.104e-05, 1.0928e-05, 1.0825e-05, 
    1.0729e-05, 1.0631e-05, 1.0535e-05, 1.0437e-05, 1.0335e-05, 1.0217e-05, 
    1.0099e-05, 9.971e-06, 9.832e-06, 9.68e-06, 9.532e-06, 9.39e-06, 
    9.255e-06, 9.144e-06, 9.044e-06, 8.946e-06, 8.852e-06, 8.759e-06, 
    8.671e-06, 8.598e-06, 8.537e-06, 8.474e-06, 8.418e-06, 8.342e-06, 
    8.244e-06, 8.131e-06, 8.012e-06, 7.915e-06, 7.828e-06, 7.757e-06, 
    7.7e-06, 7.656e-06, 7.64e-06, 7.648e-06, 7.681e-06, 7.732e-06, 7.794e-06, 
    7.863e-06, 7.938e-06, 8.033e-06, 8.155e-06, 8.264e-06, 8.383e-06, 
    8.555e-06, 8.771e-06, 9.012e-06, 9.214e-06, 9.382e-06, 9.505e-06, 
    9.608e-06, 9.638e-06, 9.612e-06, 9.54e-06, 9.42e-06, 9.268e-06, 9.09e-06, 
    8.908e-06, 8.713e-06, 8.524e-06, 8.352e-06, 8.201e-06, 8.057e-06, 
    7.927e-06, 7.806e-06, 7.693e-06, 7.613e-06, 7.566e-06, 7.533e-06, 
    7.522e-06, 7.506e-06, 7.494e-06, 7.48e-06, 7.476e-06, 7.482e-06, 
    7.463e-06, 7.418e-06, 7.331e-06, 7.201e-06, 7.044e-06, 6.869e-06, 
    6.687e-06, 6.5e-06, 6.31e-06, 6.11e-06, 5.909e-06, 5.71e-06, 5.527e-06, 
    5.355e-06, 5.199e-06, 5.068e-06, 4.958e-06, 4.861e-06, 4.773e-06, 
    4.697e-06, 4.633e-06, 4.576e-06, 4.521e-06, 4.466e-06, 4.407e-06, 
    4.35e-06, 4.296e-06, 4.24e-06, 4.194e-06, 4.151e-06, 4.128e-06, 
    4.143e-06, 4.21e-06, 4.342e-06, 4.533e-06, 4.788e-06, 5.039e-06, 
    5.281e-06, 5.509e-06, 5.692e-06, 5.865e-06, 6.039e-06, 6.182e-06, 
    6.289e-06, 6.342e-06, 6.35e-06, 6.263e-06, 6.133e-06, 5.947e-06, 
    5.683e-06, 5.356e-06, 4.967e-06, 4.536e-06, 4.079e-06, 3.61e-06, 
    3.143e-06, 2.71e-06, 2.344e-06, 2.053e-06, 1.82e-06, 1.642e-06, 
    1.535e-06, 1.541e-06, 1.634e-06, 1.829e-06, 2.119e-06, 2.468e-06, 
    2.802e-06, 3.043e-06, 3.243e-06, 3.416e-06, 3.569e-06, 3.681e-06, 
    3.799e-06, 3.883e-06, 3.948e-06, 3.999e-06, 4.015e-06, 3.984e-06, 
    3.933e-06, 3.871e-06, 3.824e-06, 3.809e-06, 3.833e-06, 3.903e-06, 
    4.015e-06, 4.146e-06, 4.297e-06, 4.433e-06, 4.566e-06, 4.67e-06, 
    4.747e-06, 4.79e-06, 4.802e-06, 4.793e-06, 4.755e-06, 4.712e-06, 
    4.637e-06, 4.542e-06, 4.429e-06, 4.292e-06, 4.129e-06, 3.952e-06, 
    3.776e-06, 3.619e-06, 3.481e-06, 3.36e-06, 3.28e-06, 3.201e-06, 
    3.136e-06, 3.08e-06, 3.031e-06, 3.009e-06, 3.007e-06, 2.995e-06, 
    2.976e-06, 2.984e-06, 3.02e-06, 3.054e-06, 3.033e-06, 2.965e-06, 
    2.863e-06, 2.763e-06, 2.696e-06, 2.671e-06, 2.693e-06, 2.742e-06, 
    2.808e-06, 2.882e-06, 2.975e-06, 3.095e-06, 3.25e-06, 3.445e-06, 
    3.648e-06, 3.841e-06, 4.033e-06, 4.212e-06, 4.361e-06, 4.461e-06, 
    4.514e-06, 4.521e-06, 4.474e-06, 4.379e-06, 4.273e-06, 4.165e-06, 
    4.054e-06, 3.955e-06, 3.873e-06, 3.796e-06, 3.695e-06, 3.594e-06, 
    3.499e-06, 3.409e-06, 3.32e-06, 3.258e-06, 3.204e-06, 3.125e-06, 
    3.029e-06, 2.911e-06, 2.79e-06, 2.665e-06, 2.558e-06, 2.464e-06, 
    2.373e-06, 2.299e-06, 2.252e-06, 2.226e-06, 2.223e-06, 2.246e-06, 
    2.296e-06, 2.352e-06, 2.416e-06, 2.474e-06, 2.516e-06, 2.553e-06, 
    2.596e-06, 2.627e-06, 2.7e-06, 2.849e-06, 3.046e-06, 3.296e-06, 
    3.556e-06, 3.817e-06, 4.008e-06, 4.103e-06, 4.08e-06, 4.015e-06, 
    3.906e-06, 3.754e-06, 3.578e-06, 3.372e-06, 3.145e-06, 2.91e-06, 
    2.692e-06, 2.501e-06, 2.341e-06, 2.21e-06, 2.119e-06, 2.048e-06, 
    1.988e-06, 1.95e-06, 1.931e-06, 1.911e-06, 1.879e-06, 1.857e-06, 
    1.843e-06, 1.823e-06, 1.804e-06, 1.787e-06, 1.77e-06, 1.751e-06, 
    1.719e-06, 1.693e-06, 1.682e-06, 1.679e-06, 1.687e-06, 1.699e-06, 
    1.74e-06, 1.803e-06, 1.889e-06, 1.981e-06, 2.083e-06, 2.174e-06, 
    2.247e-06, 2.327e-06, 2.417e-06, 2.484e-06, 2.546e-06, 2.613e-06, 
    2.662e-06, 2.702e-06, 2.734e-06, 2.769e-06, 2.807e-06, 2.849e-06, 
    2.891e-06, 2.931e-06, 2.96e-06, 2.962e-06, 2.939e-06, 2.893e-06, 
    2.831e-06, 2.749e-06, 2.657e-06, 2.56e-06, 2.442e-06, 2.325e-06, 
    2.204e-06, 2.083e-06, 1.966e-06, 1.854e-06, 1.754e-06, 1.669e-06, 
    1.6e-06, 1.545e-06, 1.505e-06, 1.476e-06, 1.455e-06, 1.445e-06, 
    1.424e-06, 1.39e-06, 1.336e-06, 1.262e-06, 1.167e-06, 1.071e-06, 
    9.75e-07, 8.91e-07, 8.18e-07, 7.64e-07, 7.35e-07, 7.29e-07, 7.34e-07, 
    7.48e-07, 7.66e-07, 7.92e-07, 8.34e-07, 8.84e-07, 9.25e-07, 9.4e-07, 
    9.28e-07, 9e-07, 8.6e-07, 8.18e-07, 7.79e-07, 7.53e-07, 7.33e-07, 
    7.14e-07, 6.96e-07, 6.77e-07, 6.67e-07, 6.66e-07, 6.61e-07, 6.58e-07, 
    6.66e-07, 6.88e-07, 7.21e-07, 7.65e-07, 8.15e-07, 8.67e-07, 9.21e-07, 
    9.87e-07, 1.086e-06, 1.224e-06, 1.378e-06, 1.525e-06, 1.663e-06, 
    1.762e-06, 1.859e-06, 1.943e-06, 2.009e-06, 2.047e-06, 2.052e-06, 
    2.012e-06, 1.937e-06, 1.819e-06, 1.677e-06, 1.522e-06, 1.361e-06, 
    1.202e-06, 1.053e-06, 9.19e-07, 7.9e-07, 6.79e-07, 5.93e-07, 5.28e-07, 
    4.99e-07, 4.83e-07, 4.68e-07, 4.43e-07, 4.02e-07, 3.56e-07, 3e-07, 
    2.35e-07, 1.84e-07, 1.53e-07, 1.38e-07, 1.53e-07, 1.74e-07, 1.99e-07, 
    2.22e-07, 2.27e-07, 2.27e-07, 2.11e-07, 1.99e-07, 1.86e-07, 1.57e-07, 
    1.3e-07, 7.7e-08, -8e-09, -1.13e-07, -2.38e-07, -3.8e-07, -5.04e-07, 
    -5.87e-07, -6.25e-07, -5.5e-07, -4.12e-07, -1.99e-07, 4.1e-08, 2.76e-07, 
    6e-07, 9.24e-07, 1.16e-06, 1.393e-06, 1.599e-06, 1.834e-06, 2.074e-06, 
    2.218e-06, 2.259e-06, 2.214e-06, 2.11e-06, 1.987e-06, 1.888e-06, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, 0.0021696, 0.0021573, 0.0021454, 
    0.0021335, 0.0021214, 0.0021092, 0.0020971, 0.0020854, 0.0020741, 
    0.002063, 0.0020521, 0.0020412, 0.0020307, 0.0020203, 0.0020099, 
    0.0019995, 0.0019901, 0.0019804, 0.0019709, 0.0019621, 0.0019529, 
    0.0019446, 0.0019365, 0.0019288, 0.0019218, 0.0019149, 0.0019084, 
    0.0019028, 0.0018967, 0.0018919, 0.0018871, 0.0018827, 0.0018789, 
    0.0018763, 0.0018732, 0.0018691, 0.0018637, 0.001858, 0.0018513, 
    0.0018435, 0.0018348, 0.0018258, 0.001816, 0.0018054, 0.0017945, 
    0.0017833, 0.0017717, 0.0017598, 0.001748, 0.0017363, 0.0017246, 
    0.0017131, 0.0017016, 0.0016906, 0.0016793, 0.0016683, 0.0016574, 
    0.0016469, 0.0016364, 0.0016259, 0.0016155, 0.0016053, 0.0015953, 
    0.0015853, 0.0015754, 0.0015655, 0.0015556, 0.0015458, 0.0015363, 
    0.0015269, 0.0015173, 0.0015078, 0.0014986, 0.0014894, 0.0014802, 
    0.0014712, 0.0014621, 0.0014529, 0.0014439, 0.0014348, 0.0014258, 
    0.0014169, 0.0014082, 0.0013996, 0.0013911, 0.0013828, 0.0013744, 
    0.0013665, 0.0013586, 0.0013508, 0.0013434, 0.0013362, 0.0013292, 
    0.001322, 0.0013152, 0.0013085, 0.0013019, 0.0012956, 0.0012893, 
    0.0012832, 0.001277, 0.001271, 0.0012652, 0.0012595, 0.0012539, 
    0.0012483, 0.0012426, 0.0012369, 0.0012307, 0.0012242, 0.0012176, 
    0.0012111, 0.0012042, 0.0011971, 0.00119, 0.001183, 0.0011759, 0.0011684, 
    0.0011609, 0.0011533, 0.0011452, 0.0011372, 0.0011292, 0.0011211, 
    0.001113, 0.0011047, 0.0010966, 0.0010886, 0.0010806, 0.001073, 
    0.0010656, 0.0010581, 0.001051, 0.001044, 0.0010371, 0.0010305, 
    0.0010242, 0.0010178, 0.0010116, 0.0010057, 0.00099995, 0.0009944, 
    0.00098904, 0.00098375, 0.00097859, 0.00097346, 0.00096835, 0.0009633, 
    0.0009582, 0.00095317, 0.00094811, 0.00094303, 0.00093786, 0.00093253, 
    0.00092711, 0.0009216, 0.00091593, 0.00091006, 0.00090409, 0.00089794, 
    0.0008916, 0.00088503, 0.00087825, 0.00087138, 0.00086437, 0.00085731, 
    0.00085019, 0.00084312, 0.00083595, 0.00082885, 0.00082148, 0.00081415, 
    0.00080699, 0.00079992, 0.00079284, 0.00078585, 0.00077893, 0.00077234, 
    0.000766, 0.00075973, 0.00075371, 0.00074774, 0.00074182, 0.00073604, 
    0.00073031, 0.00072466, 0.00071909, 0.00071351, 0.00070805, 0.00070259, 
    0.00069721, 0.00069202, 0.00068692, 0.00068183, 0.00067677, 0.00067184, 
    0.00066691, 0.00066199, 0.00065709, 0.00065221, 0.00064737, 0.0006426, 
    0.00063792, 0.00063329, 0.0006287, 0.00062413, 0.00061965, 0.00061522, 
    0.00061077, 0.00060635, 0.00060205, 0.00059786, 0.0005938, 0.00058971, 
    0.00058566, 0.00058168, 0.00057777, 0.00057394, 0.00057019, 0.00056655, 
    0.00056301, 0.00055949, 0.00055601, 0.00055251, 0.000549, 0.0005454, 
    0.0005418, 0.00053824, 0.00053468, 0.00053111, 0.00052756, 0.00052397, 
    0.00052042, 0.00051685, 0.00051326, 0.00050969, 0.0005061, 0.00050249, 
    0.0004989, 0.00049533, 0.00049175, 0.00048818, 0.00048464, 0.00048113, 
    0.00047758, 0.00047398, 0.00047036, 0.00046677, 0.00046319, 0.00045964, 
    0.00045615, 0.00045263, 0.00044912, 0.00044559, 0.00044206, 0.00043854, 
    0.0004351, 0.00043163, 0.00042814, 0.00042467, 0.00042115, 0.00041764, 
    0.00041418, 0.00041069, 0.00040723, 0.00040376, 0.00040036, 0.00039703, 
    0.00039372, 0.00039048, 0.00038732, 0.00038424, 0.0003812, 0.00037819, 
    0.00037517, 0.00037217, 0.00036926, 0.00036638, 0.0003635, 0.00036068, 
    0.0003579, 0.00035516, 0.00035247, 0.00034983, 0.00034721, 0.0003446, 
    0.00034198, 0.00033937, 0.00033675, 0.00033412, 0.00033152, 0.00032893, 
    0.00032637, 0.00032382, 0.00032128, 0.00031877, 0.00031628, 0.00031382, 
    0.00031139, 0.00030899, 0.00030661, 0.00030425, 0.00030191, 0.00029957, 
    0.00029722, 0.00029491, 0.0002926, 0.00029028, 0.00028794, 0.00028561, 
    0.00028326, 0.00028097, 0.00027875, 0.00027654, 0.00027434, 0.00027214, 
    0.00026995, 0.00026779, 0.0002656, 0.00026343, 0.00026132, 0.0002592, 
    0.00025711, 0.00025508, 0.00025301, 0.00025092, 0.0002488, 0.00024663, 
    0.00024448, 0.00024231, 0.00024014, 0.00023799, 0.00023591, 0.00023387, 
    0.00023183, 0.00022982, 0.00022778, 0.00022574, 0.00022371, 0.00022167, 
    0.00021966, 0.0002177, 0.00021578, 0.0002139, 0.00021208, 0.00021031, 
    0.00020856, 0.00020687, 0.00020522, 0.0002036, 0.00020202, 0.00020048, 
    0.00019896, 0.00019745, 0.00019594, 0.00019443, 0.00019292, 0.00019142, 
    0.00018992, 0.00018841, 0.00018692, 0.00018544, 0.00018399, 0.00018255, 
    0.00018111, 0.00017966, 0.00017822, 0.00017677, 0.00017532, 0.00017389, 
    0.00017244, 0.00017102, 0.00016964, 0.00016828, 0.00016693, 0.0001656, 
    0.00016428, 0.00016299, 0.00016171, 0.00016044, 0.0001592, 0.00015798, 
    0.00015677, 0.00015559, 0.00015442, 0.00015325, 0.00015208, 0.00015091, 
    0.00014973, 0.00014856, 0.0001474, 0.00014624, 0.00014508, 0.00014393, 
    0.00014279, 0.00014164, 0.0001405, 0.00013936, 0.00013821, 0.00013711, 
    0.00013602, 0.00013494, 0.00013388, 0.00013284, 0.00013179, 0.00013075, 
    0.00012973, 0.0001287, 0.00012765, 0.00012661, 0.00012556, 0.00012454, 
    0.00012352, 0.00012252, 0.00012153, 0.00012053, 0.00011954, 0.00011853, 
    0.00011753, 0.00011652, 0.00011551, 0.00011449, 0.00011347, 0.00011246, 
    0.00011145, 0.00011045, 0.00010945, 0.00010844, 0.00010744, 0.00010644, 
    0.00010545, 0.00010446, 0.00010347, 0.0001025, 0.00010154, 0.00010058, 
    9.9631e-05, 9.8686e-05, 9.7742e-05, 9.6814e-05, 9.5899e-05, 9.501e-05, 
    9.4148e-05, 9.3298e-05, 9.2462e-05, 9.1631e-05, 9.0856e-05, 9.0102e-05, 
    8.933e-05, 8.8552e-05, 8.7777e-05, 8.7006e-05, 8.6229e-05, 8.5462e-05, 
    8.4724e-05, 8.3997e-05, 8.3237e-05, 8.2457e-05, 8.1649e-05, 8.0825e-05, 
    8.001e-05, 7.9192e-05, 7.8386e-05, 7.7583e-05, 7.6781e-05, 7.5974e-05, 
    7.5176e-05, 7.4386e-05, 7.3609e-05, 7.2852e-05, 7.2123e-05, 7.1421e-05, 
    7.0745e-05, 7.0108e-05, 6.9496e-05, 6.8908e-05, 6.8338e-05, 6.7786e-05, 
    6.7264e-05, 6.6766e-05, 6.6283e-05, 6.5818e-05, 6.536e-05, 6.4899e-05, 
    6.4426e-05, 6.3955e-05, 6.3464e-05, 6.2965e-05, 6.2465e-05, 6.1967e-05, 
    6.1457e-05, 6.0941e-05, 6.0417e-05, 5.9882e-05, 5.9339e-05, 5.8783e-05, 
    5.8223e-05, 5.7679e-05, 5.7124e-05, 5.6564e-05, 5.6016e-05, 5.5503e-05, 
    5.4996e-05, 5.4532e-05, 5.4056e-05, 5.3599e-05, 5.3114e-05, 5.2668e-05, 
    5.2295e-05, 5.191e-05, 5.1541e-05, 5.118e-05, 5.0801e-05, 5.0415e-05, 
    5.0034e-05, 4.966e-05, 4.9297e-05, 4.8943e-05, 4.8587e-05, 4.8225e-05, 
    4.7859e-05, 4.7498e-05, 4.7138e-05, 4.6792e-05, 4.6447e-05, 4.6107e-05, 
    4.5761e-05, 4.5422e-05, 4.5084e-05, 4.4741e-05, 4.4395e-05, 4.4057e-05, 
    4.371e-05, 4.3365e-05, 4.3014e-05, 4.2656e-05, 4.2294e-05, 4.1951e-05, 
    4.1609e-05, 4.1261e-05, 4.0908e-05, 4.0552e-05, 4.0199e-05, 3.985e-05, 
    3.951e-05, 3.9165e-05, 3.8816e-05, 3.8469e-05, 3.8131e-05, 3.7808e-05, 
    3.7498e-05, 3.7207e-05, 3.6917e-05, 3.6625e-05, 3.6328e-05, 3.6027e-05, 
    3.5725e-05, 3.5422e-05, 3.5118e-05, 3.4811e-05, 3.4513e-05, 3.4212e-05, 
    3.3914e-05, 3.3615e-05, 3.331e-05, 3.3018e-05, 3.2761e-05, 3.254e-05, 
    3.2336e-05, 3.2143e-05, 3.1954e-05, 3.1765e-05, 3.1569e-05, 3.1367e-05, 
    3.116e-05, 3.0945e-05, 3.0717e-05, 3.047e-05, 3.0205e-05, 2.9928e-05, 
    2.9638e-05, 2.9347e-05, 2.9063e-05, 2.8788e-05, 2.8522e-05, 2.8262e-05, 
    2.8015e-05, 2.7783e-05, 2.7554e-05, 2.7329e-05, 2.7109e-05, 2.6894e-05, 
    2.668e-05, 2.6473e-05, 2.6284e-05, 2.6093e-05, 2.5896e-05, 2.5689e-05, 
    2.5518e-05, 2.5369e-05, 2.5224e-05, 2.5096e-05, 2.5005e-05, 2.4945e-05, 
    2.489e-05, 2.4849e-05, 2.4793e-05, 2.4748e-05, 2.4729e-05, 2.4658e-05, 
    2.4577e-05, 2.4489e-05, 2.4339e-05, 2.4139e-05, 2.3847e-05, 2.3458e-05, 
    2.2975e-05, 2.2419e-05, 2.1803e-05, 2.1151e-05, 2.0492e-05, 1.9852e-05, 
    1.9248e-05, 1.8704e-05, 1.8245e-05, 1.7891e-05, 1.7642e-05, 1.7519e-05, 
    1.7535e-05, 1.7648e-05, 1.7887e-05, 1.8239e-05, 1.8661e-05, 1.912e-05, 
    1.9594e-05, 2.0014e-05, 2.0309e-05, 2.0484e-05, 2.0523e-05, 2.0516e-05, 
    2.045e-05, 2.0319e-05, 2.0143e-05, 1.9918e-05, 1.9672e-05, 1.9428e-05, 
    1.9191e-05, 1.8978e-05, 1.8798e-05, 1.8641e-05, 1.8529e-05, 1.8457e-05, 
    1.8411e-05, 1.8412e-05, 1.8448e-05, 1.8508e-05, 1.8571e-05, 1.8608e-05, 
    1.8602e-05, 1.8575e-05, 1.8491e-05, 1.8357e-05, 1.818e-05, 1.7966e-05, 
    1.7712e-05, 1.7408e-05, 1.706e-05, 1.6678e-05, 1.6279e-05, 1.5889e-05, 
    1.5526e-05, 1.5194e-05, 1.4893e-05, 1.4627e-05, 1.4394e-05, 1.4201e-05, 
    1.4057e-05, 1.396e-05, 1.3916e-05, 1.3872e-05, 1.3848e-05, 1.3828e-05, 
    1.381e-05, 1.3786e-05, 1.3756e-05, 1.3734e-05, 1.3715e-05, 1.3697e-05, 
    1.3661e-05, 1.3607e-05, 1.3547e-05, 1.3491e-05, 1.3441e-05, 1.3389e-05, 
    1.3343e-05, 1.33e-05, 1.3257e-05, 1.3225e-05, 1.3192e-05, 1.3161e-05, 
    1.3136e-05, 1.3096e-05, 1.305e-05, 1.2999e-05, 1.2938e-05, 1.2867e-05, 
    1.2771e-05, 1.267e-05, 1.2584e-05, 1.2524e-05, 1.248e-05, 1.2439e-05, 
    1.2376e-05, 1.2271e-05, 1.2134e-05, 1.1979e-05, 1.1808e-05, 1.1633e-05, 
    1.1461e-05, 1.1306e-05, 1.1165e-05, 1.104e-05, 1.0928e-05, 1.0825e-05, 
    1.0729e-05, 1.0631e-05, 1.0535e-05, 1.0437e-05, 1.0335e-05, 1.0217e-05, 
    1.0099e-05, 9.971e-06, 9.832e-06, 9.68e-06, 9.532e-06, 9.39e-06, 
    9.255e-06, 9.144e-06, 9.044e-06, 8.946e-06, 8.852e-06, 8.759e-06, 
    8.671e-06, 8.598e-06, 8.537e-06, 8.474e-06, 8.418e-06, 8.342e-06, 
    8.244e-06, 8.131e-06, 8.012e-06, 7.915e-06, 7.828e-06, 7.757e-06, 
    7.7e-06, 7.656e-06, 7.64e-06, 7.648e-06, 7.681e-06, 7.732e-06, 7.794e-06, 
    7.863e-06, 7.938e-06, 8.033e-06, 8.155e-06, 8.264e-06, 8.383e-06, 
    8.555e-06, 8.771e-06, 9.012e-06, 9.214e-06, 9.382e-06, 9.505e-06, 
    9.608e-06, 9.638e-06, 9.612e-06, 9.54e-06, 9.42e-06, 9.268e-06, 9.09e-06, 
    8.908e-06, 8.713e-06, 8.524e-06, 8.352e-06, 8.201e-06, 8.057e-06, 
    7.927e-06, 7.806e-06, 7.693e-06, 7.613e-06, 7.566e-06, 7.533e-06, 
    7.522e-06, 7.506e-06, 7.494e-06, 7.48e-06, 7.476e-06, 7.482e-06, 
    7.463e-06, 7.418e-06, 7.331e-06, 7.201e-06, 7.044e-06, 6.869e-06, 
    6.687e-06, 6.5e-06, 6.31e-06, 6.11e-06, 5.909e-06, 5.71e-06, 5.527e-06, 
    5.355e-06, 5.199e-06, 5.068e-06, 4.958e-06, 4.861e-06, 4.773e-06, 
    4.697e-06, 4.633e-06, 4.576e-06, 4.521e-06, 4.466e-06, 4.407e-06, 
    4.35e-06, 4.296e-06, 4.24e-06, 4.194e-06, 4.151e-06, 4.128e-06, 
    4.143e-06, 4.21e-06, 4.342e-06, 4.533e-06, 4.788e-06, 5.039e-06, 
    5.281e-06, 5.509e-06, 5.692e-06, 5.865e-06, 6.039e-06, 6.182e-06, 
    6.289e-06, 6.342e-06, 6.35e-06, 6.263e-06, 6.133e-06, 5.947e-06, 
    5.683e-06, 5.356e-06, 4.967e-06, 4.536e-06, 4.079e-06, 3.61e-06, 
    3.143e-06, 2.71e-06, 2.344e-06, 2.053e-06, 1.82e-06, 1.642e-06, 
    1.535e-06, 1.541e-06, 1.634e-06, 1.829e-06, 2.119e-06, 2.468e-06, 
    2.802e-06, 3.043e-06, 3.243e-06, 3.416e-06, 3.569e-06, 3.681e-06, 
    3.799e-06, 3.883e-06, 3.948e-06, 3.999e-06, 4.015e-06, 3.984e-06, 
    3.933e-06, 3.871e-06, 3.824e-06, 3.809e-06, 3.833e-06, 3.903e-06, 
    4.015e-06, 4.146e-06, 4.297e-06, 4.433e-06, 4.566e-06, 4.67e-06, 
    4.747e-06, 4.79e-06, 4.802e-06, 4.793e-06, 4.755e-06, 4.712e-06, 
    4.637e-06, 4.542e-06, 4.429e-06, 4.292e-06, 4.129e-06, 3.952e-06, 
    3.776e-06, 3.619e-06, 3.481e-06, 3.36e-06, 3.28e-06, 3.201e-06, 
    3.136e-06, 3.08e-06, 3.031e-06, 3.009e-06, 3.007e-06, 2.995e-06, 
    2.976e-06, 2.984e-06, 3.02e-06, 3.054e-06, 3.033e-06, 2.965e-06, 
    2.863e-06, 2.763e-06, 2.696e-06, 2.671e-06, 2.693e-06, 2.742e-06, 
    2.808e-06, 2.882e-06, 2.975e-06, 3.095e-06, 3.25e-06, 3.445e-06, 
    3.648e-06, 3.841e-06, 4.033e-06, 4.212e-06, 4.361e-06, 4.461e-06, 
    4.514e-06, 4.521e-06, 4.474e-06, 4.379e-06, 4.273e-06, 4.165e-06, 
    4.054e-06, 3.955e-06, 3.873e-06, 3.796e-06, 3.695e-06, 3.594e-06, 
    3.499e-06, 3.409e-06, 3.32e-06, 3.258e-06, 3.204e-06, 3.125e-06, 
    3.029e-06, 2.911e-06, 2.79e-06, 2.665e-06, 2.558e-06, 2.464e-06, 
    2.373e-06, 2.299e-06, 2.252e-06, 2.226e-06, 2.223e-06, 2.246e-06, 
    2.296e-06, 2.352e-06, 2.416e-06, 2.474e-06, 2.516e-06, 2.553e-06, 
    2.596e-06, 2.627e-06, 2.7e-06, 2.849e-06, 3.046e-06, 3.296e-06, 
    3.556e-06, 3.817e-06, 4.008e-06, 4.103e-06, 4.08e-06, 4.015e-06, 
    3.906e-06, 3.754e-06, 3.578e-06, 3.372e-06, 3.145e-06, 2.91e-06, 
    2.692e-06, 2.501e-06, 2.341e-06, 2.21e-06, 2.119e-06, 2.048e-06, 
    1.988e-06, 1.95e-06, 1.931e-06, 1.911e-06, 1.879e-06, 1.857e-06, 
    1.843e-06, 1.823e-06, 1.804e-06, 1.787e-06, 1.77e-06, 1.751e-06, 
    1.719e-06, 1.693e-06, 1.682e-06, 1.679e-06, 1.687e-06, 1.699e-06, 
    1.74e-06, 1.803e-06, 1.889e-06, 1.981e-06, 2.083e-06, 2.174e-06, 
    2.247e-06, 2.327e-06, 2.417e-06, 2.484e-06, 2.546e-06, 2.613e-06, 
    2.662e-06, 2.702e-06, 2.734e-06, 2.769e-06, 2.807e-06, 2.849e-06, 
    2.891e-06, 2.931e-06, 2.96e-06, 2.962e-06, 2.939e-06, 2.893e-06, 
    2.831e-06, 2.749e-06, 2.657e-06, 2.56e-06, 2.442e-06, 2.325e-06, 
    2.204e-06, 2.083e-06, 1.966e-06, 1.854e-06, 1.754e-06, 1.669e-06, 
    1.6e-06, 1.545e-06, 1.505e-06, 1.476e-06, 1.455e-06, 1.445e-06, 
    1.424e-06, 1.39e-06, 1.336e-06, 1.262e-06, 1.167e-06, 1.071e-06, 
    9.75e-07, 8.91e-07, 8.18e-07, 7.64e-07, 7.35e-07, 7.29e-07, 7.34e-07, 
    7.48e-07, 7.66e-07, 7.92e-07, 8.34e-07, 8.84e-07, 9.25e-07, 9.4e-07, 
    9.28e-07, 9e-07, 8.6e-07, 8.18e-07, 7.79e-07, 7.53e-07, 7.33e-07, 
    7.14e-07, 6.96e-07, 6.77e-07, 6.67e-07, 6.66e-07, 6.61e-07, 6.58e-07, 
    6.66e-07, 6.88e-07, 7.21e-07, 7.65e-07, 8.15e-07, 8.67e-07, 9.21e-07, 
    9.87e-07, 1.086e-06, 1.224e-06, 1.378e-06, 1.525e-06, 1.663e-06, 
    1.762e-06, 1.859e-06, 1.943e-06, 2.009e-06, 2.047e-06, 2.052e-06, 
    2.012e-06, 1.937e-06, 1.819e-06, 1.677e-06, 1.522e-06, 1.361e-06, 
    1.202e-06, 1.053e-06, 9.19e-07, 7.9e-07, 6.79e-07, 5.93e-07, 5.28e-07, 
    4.99e-07, 4.83e-07, 4.68e-07, 4.43e-07, 4.02e-07, 3.56e-07, 3e-07, 
    2.35e-07, 1.84e-07, 1.53e-07, 1.38e-07, 1.53e-07, 1.74e-07, 1.99e-07, 
    2.22e-07, 2.27e-07, 2.27e-07, 2.11e-07, 1.99e-07, 1.86e-07, 1.57e-07, 
    1.3e-07, 7.7e-08, -8e-09, -1.13e-07, -2.38e-07, -3.8e-07, -5.04e-07, 
    -5.87e-07, -6.25e-07, -5.5e-07, -4.12e-07, -1.99e-07, 4.1e-08, 2.76e-07, 
    6e-07, 9.24e-07, 1.16e-06, 1.393e-06, 1.599e-06, 1.834e-06, 2.074e-06, 
    2.218e-06, 2.259e-06, 2.214e-06, 2.11e-06, 1.987e-06, 1.888e-06, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L1_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_L2_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 bangle_opt_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07 ;

 alt_refrac =
  18263, 18365, 18468, 18571, 18673, 18776, 18879, 18981, 19084, 19186, 
    19289, 19391, 19494, 19596, 19698, 19800, 19902, 20004, 20106, 20207, 
    20309, 20411, 20513, 20615, 20716, 20818, 20920, 21022, 21123, 21225, 
    21327, 21428, 21530, 21631, 21733, 21834, 21936, 22037, 22139, 22240, 
    22342, 22443, 22544, 22646, 22747, 22848, 22950, 23051, 23152, 23253, 
    23354, 23455, 23556, 23658, 23759, 23860, 23961, 24062, 24163, 24264, 
    24365, 24467, 24568, 24669, 24770, 24871, 24972, 25072, 25173, 25274, 
    25375, 25476, 25576, 25677, 25778, 25879, 25979, 26080, 26181, 26281, 
    26382, 26483, 26583, 26684, 26785, 26885, 26986, 27086, 27187, 27288, 
    27388, 27489, 27589, 27690, 27790, 27891, 27991, 28092, 28192, 28293, 
    28393, 28494, 28594, 28695, 28795, 28896, 28996, 29097, 29197, 29297, 
    29398, 29498, 29599, 29699, 29799, 29900, 30000, 30100, 30201, 30301, 
    30401, 30502, 30602, 30702, 30803, 30903, 31003, 31104, 31204, 31304, 
    31404, 31505, 31605, 31705, 31806, 31906, 32006, 32106, 32207, 32307, 
    32407, 32507, 32608, 32708, 32808, 32908, 33008, 33108, 33209, 33309, 
    33409, 33509, 33609, 33710, 33810, 33910, 34010, 34110, 34210, 34310, 
    34411, 34511, 34611, 34711, 34811, 34911, 35011, 35112, 35212, 35312, 
    35412, 35512, 35612, 35712, 35812, 35912, 36012, 36113, 36213, 36313, 
    36413, 36513, 36613, 36713, 36813, 36913, 37014, 37114, 37214, 37314, 
    37414, 37514, 37614, 37714, 37814, 37914, 38014, 38114, 38214, 38314, 
    38414, 38514, 38614, 38715, 38815, 38915, 39015, 39115, 39215, 39315, 
    39415, 39515, 39615, 39715, 39815, 39915, 40015, 40115, 40215, 40315, 
    40415, 40515, 40615, 40715, 40815, 40915, 41015, 41115, 41215, 41315, 
    41415, 41515, 41615, 41715, 41815, 41915, 42015, 42115, 42215, 42315, 
    42415, 42515, 42615, 42715, 42815, 42915, 43015, 43115, 43215, 43315, 
    43415, 43515, 43615, 43715, 43815, 43915, 44015, 44115, 44215, 44315, 
    44415, 44515, 44615, 44715, 44815, 44915, 45015, 45115, 45215, 45315, 
    45415, 45515, 45615, 45714, 45814, 45914, 46014, 46114, 46214, 46314, 
    46414, 46514, 46614, 46714, 46814, 46914, 47014, 47114, 47214, 47314, 
    47414, 47514, 47614, 47714, 47814, 47914, 48014, 48114, 48214, 48314, 
    48414, 48514, 48614, 48714, 48813, 48913, 49013, 49113, 49213, 49313, 
    49413, 49513, 49613, 49713, 49813, 49913, 50013, 50113, 50213, 50313, 
    50413, 50513, 50613, 50712, 50812, 50912, 51012, 51112, 51212, 51312, 
    51412, 51512, 51612, 51712, 51812, 51912, 52012, 52112, 52212, 52312, 
    52412, 52512, 52612, 52712, 52812, 52911, 53011, 53111, 53211, 53311, 
    53411, 53511, 53611, 53711, 53811, 53911, 54011, 54111, 54211, 54311, 
    54411, 54511, 54610, 54710, 54810, 54910, 55010, 55110, 55210, 55310, 
    55410, 55510, 55610, 55710, 55810, 55910, 56010, 56110, 56210, 56310, 
    56410, 56509, 56609, 56709, 56809, 56909, 57009, 57109, 57209, 57309, 
    57409, 57509, 57609, 57709, 57809, 57909, 58009, 58108, 58208, 58308, 
    58408, 58508, 58608, 58708, 58808, 58908, 59008, 59108, 59208, 59308, 
    59408, 59508, 59608, 59708, 59808, 59907, 60007, 60107, 60207, 60307, 
    60407, 60507, 60607, 60707, 60807, 60907, 61007, 61107, 61207, 61307, 
    61406, 61506, 61606, 61706, 61806, 61906, 62006, 62106, 62206, 62306, 
    62406, 62506, 62606, 62706, 62806, 62906, 63006, 63105, 63205, 63305, 
    63405, 63505, 63605, 63705, 63805, 63905, 64005, 64105, 64205, 64305, 
    64405, 64505, 64604, 64704, 64804, 64904, 65004, 65104, 65204, 65304, 
    65404, 65504, 65604, 65704, 65804, 65904, 66004, 66104, 66204, 66303, 
    66403, 66503, 66603, 66703, 66803, 66903, 67003, 67103, 67203, 67303, 
    67403, 67503, 67603, 67702, 67802, 67902, 68002, 68102, 68202, 68302, 
    68402, 68502, 68602, 68702, 68802, 68902, 69002, 69102, 69202, 69302, 
    69401, 69501, 69601, 69701, 69801, 69901, 70001, 70101, 70201, 70301, 
    70401, 70501, 70601, 70701, 70800, 70900, 71000, 71100, 71200, 71300, 
    71400, 71500, 71600, 71700, 71800, 71900, 72000, 72100, 72200, 72300, 
    72399, 72499, 72599, 72699, 72799, 72899, 72999, 73099, 73199, 73299, 
    73399, 73499, 73599, 73699, 73798, 73898, 73998, 74098, 74198, 74298, 
    74398, 74498, 74598, 74698, 74798, 74898, 74998, 75098, 75198, 75298, 
    75398, 75497, 75597, 75697, 75797, 75897, 75997, 76097, 76197, 76297, 
    76397, 76497, 76597, 76697, 76796, 76896, 76996, 77096, 77196, 77296, 
    77396, 77496, 77596, 77696, 77796, 77896, 77996, 78096, 78196, 78296, 
    78396, 78495, 78595, 78695, 78795, 78895, 78995, 79095, 79195, 79295, 
    79395, 79495, 79595, 79695, 79794, 79894, 79994, 80094, 80194, 80294, 
    80394, 80494, 80594, 80694, 80794, 80894, 80994, 81094, 81194, 81294, 
    81394, 81493, 81593, 81693, 81793, 81893, 81993, 82093, 82193, 82293, 
    82393, 82493, 82593, 82693, 82792, 82892, 82992, 83092, 83192, 83292, 
    83392, 83492, 83592, 83692, 83792, 83892, 83992, 84092, 84192, 84292, 
    84392, 84491, 84591, 84691, 84791, 84891, 84991, 85091, 85191, 85291, 
    85391, 85491, 85591, 85691, 85790, 85890, 85990, 86090, 86190, 86290, 
    86390, 86490, 86590, 86690, 86790, 86890, 86990, 87090, 87190, 87290, 
    87390, 87489, 87589, 87689, 87789, 87889, 87989, 88089, 88189, 88289, 
    88389, 88489, 88589, 88689, 88788, 88888, 88988, 89088, 89188, 89288, 
    89388, 89488, 89588, 89688, 89788, 89888, 89988, 90088, 90188, 90288, 
    90388, 90487, 90587, 90687, 90787, 90887, 90987, 91087, 91187, 91287, 
    91387, 91487, 91587, 91687, 91786, 91886, 91986, 92086, 92186, 92286, 
    92386, 92486, 92586, 92686, 92786, 92886, 92986, 93086, 93186, 93286, 
    93386, 93485, 93585, 93685, 93785, 93885, 93985, 94085, 94185, 94285, 
    94385, 94485, 94585, 94685, 94784, 94884, 94984, 95084, 95184, 95284, 
    95384, 95484, 95584, 95684, 95784, 95884, 95984, 96084, 96184, 96284, 
    96383, 96483, 96583, 96683, 96783, 96883, 96983, 97083, 97183, 97283, 
    97383, 97483, 97583, 97683, 97782, 97882, 97982, 98082, 98182, 98282, 
    98382, 98482, 98582, 98682, 98782, 98882, 98982, 99082, 99182, 99282, 
    99381, 99481, 99581, 99681, 99781, 99881, 99981,
  18263, 18365, 18468, 18571, 18673, 18776, 18879, 18981, 19084, 19186, 
    19289, 19391, 19494, 19596, 19698, 19800, 19902, 20004, 20106, 20207, 
    20309, 20411, 20513, 20615, 20716, 20818, 20920, 21022, 21123, 21225, 
    21327, 21428, 21530, 21631, 21733, 21834, 21936, 22037, 22139, 22240, 
    22342, 22443, 22544, 22646, 22747, 22848, 22950, 23051, 23152, 23253, 
    23354, 23455, 23556, 23658, 23759, 23860, 23961, 24062, 24163, 24264, 
    24365, 24467, 24568, 24669, 24770, 24871, 24972, 25072, 25173, 25274, 
    25375, 25476, 25576, 25677, 25778, 25879, 25979, 26080, 26181, 26281, 
    26382, 26483, 26583, 26684, 26785, 26885, 26986, 27086, 27187, 27288, 
    27388, 27489, 27589, 27690, 27790, 27891, 27991, 28092, 28192, 28293, 
    28393, 28494, 28594, 28695, 28795, 28896, 28996, 29097, 29197, 29297, 
    29398, 29498, 29599, 29699, 29799, 29900, 30000, 30100, 30201, 30301, 
    30401, 30502, 30602, 30702, 30803, 30903, 31003, 31104, 31204, 31304, 
    31404, 31505, 31605, 31705, 31806, 31906, 32006, 32106, 32207, 32307, 
    32407, 32507, 32608, 32708, 32808, 32908, 33008, 33108, 33209, 33309, 
    33409, 33509, 33609, 33710, 33810, 33910, 34010, 34110, 34210, 34310, 
    34411, 34511, 34611, 34711, 34811, 34911, 35011, 35112, 35212, 35312, 
    35412, 35512, 35612, 35712, 35812, 35912, 36012, 36113, 36213, 36313, 
    36413, 36513, 36613, 36713, 36813, 36913, 37014, 37114, 37214, 37314, 
    37414, 37514, 37614, 37714, 37814, 37914, 38014, 38114, 38214, 38314, 
    38414, 38514, 38614, 38715, 38815, 38915, 39015, 39115, 39215, 39315, 
    39415, 39515, 39615, 39715, 39815, 39915, 40015, 40115, 40215, 40315, 
    40415, 40515, 40615, 40715, 40815, 40915, 41015, 41115, 41215, 41315, 
    41415, 41515, 41615, 41715, 41815, 41915, 42015, 42115, 42215, 42315, 
    42415, 42515, 42615, 42715, 42815, 42915, 43015, 43115, 43215, 43315, 
    43415, 43515, 43615, 43715, 43815, 43915, 44015, 44115, 44215, 44315, 
    44415, 44515, 44615, 44715, 44815, 44915, 45015, 45115, 45215, 45315, 
    45415, 45515, 45615, 45714, 45814, 45914, 46014, 46114, 46214, 46314, 
    46414, 46514, 46614, 46714, 46814, 46914, 47014, 47114, 47214, 47314, 
    47414, 47514, 47614, 47714, 47814, 47914, 48014, 48114, 48214, 48314, 
    48414, 48514, 48614, 48714, 48813, 48913, 49013, 49113, 49213, 49313, 
    49413, 49513, 49613, 49713, 49813, 49913, 50013, 50113, 50213, 50313, 
    50413, 50513, 50613, 50712, 50812, 50912, 51012, 51112, 51212, 51312, 
    51412, 51512, 51612, 51712, 51812, 51912, 52012, 52112, 52212, 52312, 
    52412, 52512, 52612, 52712, 52812, 52911, 53011, 53111, 53211, 53311, 
    53411, 53511, 53611, 53711, 53811, 53911, 54011, 54111, 54211, 54311, 
    54411, 54511, 54610, 54710, 54810, 54910, 55010, 55110, 55210, 55310, 
    55410, 55510, 55610, 55710, 55810, 55910, 56010, 56110, 56210, 56310, 
    56410, 56509, 56609, 56709, 56809, 56909, 57009, 57109, 57209, 57309, 
    57409, 57509, 57609, 57709, 57809, 57909, 58009, 58108, 58208, 58308, 
    58408, 58508, 58608, 58708, 58808, 58908, 59008, 59108, 59208, 59308, 
    59408, 59508, 59608, 59708, 59808, 59907, 60007, 60107, 60207, 60307, 
    60407, 60507, 60607, 60707, 60807, 60907, 61007, 61107, 61207, 61307, 
    61406, 61506, 61606, 61706, 61806, 61906, 62006, 62106, 62206, 62306, 
    62406, 62506, 62606, 62706, 62806, 62906, 63006, 63105, 63205, 63305, 
    63405, 63505, 63605, 63705, 63805, 63905, 64005, 64105, 64205, 64305, 
    64405, 64505, 64604, 64704, 64804, 64904, 65004, 65104, 65204, 65304, 
    65404, 65504, 65604, 65704, 65804, 65904, 66004, 66104, 66204, 66303, 
    66403, 66503, 66603, 66703, 66803, 66903, 67003, 67103, 67203, 67303, 
    67403, 67503, 67603, 67702, 67802, 67902, 68002, 68102, 68202, 68302, 
    68402, 68502, 68602, 68702, 68802, 68902, 69002, 69102, 69202, 69302, 
    69401, 69501, 69601, 69701, 69801, 69901, 70001, 70101, 70201, 70301, 
    70401, 70501, 70601, 70701, 70800, 70900, 71000, 71100, 71200, 71300, 
    71400, 71500, 71600, 71700, 71800, 71900, 72000, 72100, 72200, 72300, 
    72399, 72499, 72599, 72699, 72799, 72899, 72999, 73099, 73199, 73299, 
    73399, 73499, 73599, 73699, 73798, 73898, 73998, 74098, 74198, 74298, 
    74398, 74498, 74598, 74698, 74798, 74898, 74998, 75098, 75198, 75298, 
    75398, 75497, 75597, 75697, 75797, 75897, 75997, 76097, 76197, 76297, 
    76397, 76497, 76597, 76697, 76796, 76896, 76996, 77096, 77196, 77296, 
    77396, 77496, 77596, 77696, 77796, 77896, 77996, 78096, 78196, 78296, 
    78396, 78495, 78595, 78695, 78795, 78895, 78995, 79095, 79195, 79295, 
    79395, 79495, 79595, 79695, 79794, 79894, 79994, 80094, 80194, 80294, 
    80394, 80494, 80594, 80694, 80794, 80894, 80994, 81094, 81194, 81294, 
    81394, 81493, 81593, 81693, 81793, 81893, 81993, 82093, 82193, 82293, 
    82393, 82493, 82593, 82693, 82792, 82892, 82992, 83092, 83192, 83292, 
    83392, 83492, 83592, 83692, 83792, 83892, 83992, 84092, 84192, 84292, 
    84392, 84491, 84591, 84691, 84791, 84891, 84991, 85091, 85191, 85291, 
    85391, 85491, 85591, 85691, 85790, 85890, 85990, 86090, 86190, 86290, 
    86390, 86490, 86590, 86690, 86790, 86890, 86990, 87090, 87190, 87290, 
    87390, 87489, 87589, 87689, 87789, 87889, 87989, 88089, 88189, 88289, 
    88389, 88489, 88589, 88689, 88788, 88888, 88988, 89088, 89188, 89288, 
    89388, 89488, 89588, 89688, 89788, 89888, 89988, 90088, 90188, 90288, 
    90388, 90487, 90587, 90687, 90787, 90887, 90987, 91087, 91187, 91287, 
    91387, 91487, 91587, 91687, 91786, 91886, 91986, 92086, 92186, 92286, 
    92386, 92486, 92586, 92686, 92786, 92886, 92986, 93086, 93186, 93286, 
    93386, 93485, 93585, 93685, 93785, 93885, 93985, 94085, 94185, 94285, 
    94385, 94485, 94585, 94685, 94784, 94884, 94984, 95084, 95184, 95284, 
    95384, 95484, 95584, 95684, 95784, 95884, 95984, 96084, 96184, 96284, 
    96383, 96483, 96583, 96683, 96783, 96883, 96983, 97083, 97183, 97283, 
    97383, 97483, 97583, 97683, 97782, 97882, 97982, 98082, 98182, 98282, 
    98382, 98482, 98582, 98682, 98782, 98882, 98982, 99082, 99182, 99282, 
    99381, 99481, 99581, 99681, 99781, 99881, 99981 ;

 geop_refrac =
  18219, 18321, 18423, 18526, 18628, 18730, 18832, 18934, 19036, 19138, 
    19240, 19342, 19443, 19545, 19646, 19748, 19849, 19950, 20052, 20153, 
    20254, 20355, 20457, 20558, 20659, 20760, 20861, 20962, 21063, 21164, 
    21265, 21366, 21467, 21568, 21669, 21770, 21871, 21971, 22072, 22173, 
    22274, 22375, 22475, 22576, 22677, 22777, 22878, 22978, 23079, 23179, 
    23280, 23380, 23481, 23581, 23681, 23782, 23882, 23983, 24083, 24184, 
    24284, 24384, 24485, 24585, 24685, 24785, 24886, 24986, 25086, 25186, 
    25286, 25386, 25486, 25586, 25686, 25786, 25886, 25986, 26086, 26186, 
    26286, 26385, 26485, 26585, 26685, 26785, 26884, 26984, 27084, 27184, 
    27283, 27383, 27483, 27583, 27682, 27782, 27882, 27982, 28081, 28181, 
    28280, 28380, 28480, 28579, 28679, 28778, 28878, 28978, 29077, 29177, 
    29276, 29376, 29475, 29575, 29674, 29774, 29873, 29973, 30072, 30171, 
    30271, 30370, 30470, 30569, 30668, 30768, 30867, 30967, 31066, 31165, 
    31265, 31364, 31463, 31563, 31662, 31761, 31861, 31960, 32059, 32158, 
    32258, 32357, 32456, 32555, 32655, 32754, 32853, 32952, 33051, 33151, 
    33250, 33349, 33448, 33547, 33646, 33746, 33845, 33944, 34043, 34142, 
    34241, 34340, 34439, 34538, 34638, 34737, 34836, 34935, 35034, 35133, 
    35232, 35331, 35430, 35529, 35628, 35727, 35826, 35925, 36024, 36123, 
    36222, 36321, 36420, 36519, 36618, 36717, 36816, 36915, 37014, 37113, 
    37212, 37311, 37410, 37509, 37608, 37707, 37805, 37904, 38003, 38102, 
    38201, 38300, 38399, 38498, 38597, 38696, 38794, 38893, 38992, 39091, 
    39190, 39289, 39387, 39486, 39585, 39684, 39783, 39881, 39980, 40079, 
    40178, 40277, 40375, 40474, 40573, 40672, 40771, 40869, 40968, 41067, 
    41166, 41264, 41363, 41462, 41561, 41659, 41758, 41857, 41956, 42054, 
    42153, 42252, 42350, 42449, 42548, 42646, 42745, 42844, 42942, 43041, 
    43140, 43238, 43337, 43436, 43534, 43633, 43732, 43830, 43929, 44028, 
    44126, 44225, 44324, 44422, 44521, 44619, 44718, 44817, 44915, 45014, 
    45112, 45211, 45310, 45408, 45507, 45605, 45704, 45802, 45901, 46000, 
    46098, 46197, 46295, 46394, 46492, 46591, 46689, 46788, 46886, 46985, 
    47084, 47182, 47281, 47379, 47478, 47576, 47675, 47773, 47872, 47970, 
    48069, 48167, 48266, 48364, 48462, 48561, 48659, 48758, 48856, 48955, 
    49053, 49152, 49250, 49349, 49447, 49545, 49644, 49742, 49841, 49939, 
    50038, 50136, 50234, 50333, 50431, 50530, 50628, 50726, 50825, 50923, 
    51022, 51120, 51218, 51317, 51415, 51513, 51612, 51710, 51809, 51907, 
    52005, 52104, 52202, 52300, 52399, 52497, 52595, 52694, 52792, 52890, 
    52989, 53087, 53185, 53283, 53382, 53480, 53578, 53677, 53775, 53873, 
    53972, 54070, 54168, 54266, 54365, 54463, 54561, 54659, 54758, 54856, 
    54954, 55052, 55151, 55249, 55347, 55445, 55544, 55642, 55740, 55838, 
    55937, 56035, 56133, 56231, 56329, 56428, 56526, 56624, 56722, 56820, 
    56919, 57017, 57115, 57213, 57311, 57409, 57508, 57606, 57704, 57802, 
    57900, 57998, 58097, 58195, 58293, 58391, 58489, 58587, 58685, 58784, 
    58882, 58980, 59078, 59176, 59274, 59372, 59470, 59568, 59666, 59765, 
    59863, 59961, 60059, 60157, 60255, 60353, 60451, 60549, 60647, 60745, 
    60843, 60941, 61040, 61138, 61236, 61334, 61432, 61530, 61628, 61726, 
    61824, 61922, 62020, 62118, 62216, 62314, 62412, 62510, 62608, 62706, 
    62804, 62902, 63000, 63098, 63196, 63294, 63392, 63490, 63588, 63686, 
    63784, 63882, 63980, 64077, 64175, 64273, 64371, 64469, 64567, 64665, 
    64763, 64861, 64959, 65057, 65155, 65253, 65351, 65448, 65546, 65644, 
    65742, 65840, 65938, 66036, 66134, 66232, 66330, 66427, 66525, 66623, 
    66721, 66819, 66917, 67015, 67112, 67210, 67308, 67406, 67504, 67602, 
    67700, 67797, 67895, 67993, 68091, 68189, 68286, 68384, 68482, 68580, 
    68678, 68775, 68873, 68971, 69069, 69167, 69264, 69362, 69460, 69558, 
    69656, 69753, 69851, 69949, 70047, 70144, 70242, 70340, 70438, 70535, 
    70633, 70731, 70829, 70926, 71024, 71122, 71219, 71317, 71415, 71513, 
    71610, 71708, 71806, 71903, 72001, 72099, 72197, 72294, 72392, 72490, 
    72587, 72685, 72783, 72880, 72978, 73076, 73173, 73271, 73369, 73466, 
    73564, 73662, 73759, 73857, 73954, 74052, 74150, 74247, 74345, 74442, 
    74540, 74638, 74735, 74833, 74931, 75028, 75126, 75223, 75321, 75419, 
    75516, 75614, 75711, 75809, 75906, 76004, 76102, 76199, 76297, 76394, 
    76492, 76589, 76687, 76784, 76882, 76979, 77077, 77175, 77272, 77370, 
    77467, 77565, 77662, 77760, 77857, 77955, 78052, 78150, 78247, 78345, 
    78442, 78540, 78637, 78735, 78832, 78930, 79027, 79124, 79222, 79319, 
    79417, 79514, 79612, 79709, 79807, 79904, 80001, 80099, 80196, 80294, 
    80391, 80489, 80586, 80683, 80781, 80878, 80976, 81073, 81170, 81268, 
    81365, 81463, 81560, 81657, 81755, 81852, 81950, 82047, 82144, 82242, 
    82339, 82436, 82534, 82631, 82728, 82826, 82923, 83020, 83118, 83215, 
    83312, 83410, 83507, 83604, 83702, 83799, 83896, 83994, 84091, 84188, 
    84286, 84383, 84480, 84577, 84675, 84772, 84869, 84967, 85064, 85161, 
    85258, 85356, 85453, 85550, 85647, 85745, 85842, 85939, 86036, 86134, 
    86231, 86328, 86425, 86523, 86620, 86717, 86814, 86911, 87009, 87106, 
    87203, 87300, 87398, 87495, 87592, 87689, 87786, 87883, 87981, 88078, 
    88175, 88272, 88369, 88466, 88564, 88661, 88758, 88855, 88952, 89049, 
    89147, 89244, 89341, 89438, 89535, 89632, 89729, 89826, 89924, 90021, 
    90118, 90215, 90312, 90409, 90506, 90603, 90700, 90797, 90895, 90992, 
    91089, 91186, 91283, 91380, 91477, 91574, 91671, 91768, 91865, 91962, 
    92059, 92156, 92253, 92351, 92448, 92545, 92642, 92739, 92836, 92933, 
    93030, 93127, 93224, 93321, 93418, 93515, 93612, 93709, 93806, 93903, 
    94000, 94097, 94194, 94291, 94388, 94485, 94581, 94678, 94775, 94872, 
    94969, 95066, 95163, 95260, 95357, 95454, 95551, 95648, 95745, 95842, 
    95939, 96036, 96132, 96229, 96326, 96423, 96520, 96617, 96714, 96811, 
    96908, 97005, 97102, 97198, 97295, 97392, 97489, 97586, 97683, 97780, 
    97876, 97973, 98070, 98167, 98264, 98361, 98458,
  18219, 18321, 18423, 18526, 18628, 18730, 18832, 18934, 19036, 19138, 
    19240, 19342, 19443, 19545, 19646, 19748, 19849, 19950, 20052, 20153, 
    20254, 20355, 20457, 20558, 20659, 20760, 20861, 20962, 21063, 21164, 
    21265, 21366, 21467, 21568, 21669, 21770, 21871, 21971, 22072, 22173, 
    22274, 22375, 22475, 22576, 22677, 22777, 22878, 22978, 23079, 23179, 
    23280, 23380, 23481, 23581, 23681, 23782, 23882, 23983, 24083, 24184, 
    24284, 24384, 24485, 24585, 24685, 24785, 24886, 24986, 25086, 25186, 
    25286, 25386, 25486, 25586, 25686, 25786, 25886, 25986, 26086, 26186, 
    26286, 26385, 26485, 26585, 26685, 26785, 26884, 26984, 27084, 27184, 
    27283, 27383, 27483, 27583, 27682, 27782, 27882, 27982, 28081, 28181, 
    28280, 28380, 28480, 28579, 28679, 28778, 28878, 28978, 29077, 29177, 
    29276, 29376, 29475, 29575, 29674, 29774, 29873, 29973, 30072, 30171, 
    30271, 30370, 30470, 30569, 30668, 30768, 30867, 30967, 31066, 31165, 
    31265, 31364, 31463, 31563, 31662, 31761, 31861, 31960, 32059, 32158, 
    32258, 32357, 32456, 32555, 32655, 32754, 32853, 32952, 33051, 33151, 
    33250, 33349, 33448, 33547, 33646, 33746, 33845, 33944, 34043, 34142, 
    34241, 34340, 34439, 34538, 34638, 34737, 34836, 34935, 35034, 35133, 
    35232, 35331, 35430, 35529, 35628, 35727, 35826, 35925, 36024, 36123, 
    36222, 36321, 36420, 36519, 36618, 36717, 36816, 36915, 37014, 37113, 
    37212, 37311, 37410, 37509, 37608, 37707, 37805, 37904, 38003, 38102, 
    38201, 38300, 38399, 38498, 38597, 38696, 38794, 38893, 38992, 39091, 
    39190, 39289, 39387, 39486, 39585, 39684, 39783, 39881, 39980, 40079, 
    40178, 40277, 40375, 40474, 40573, 40672, 40771, 40869, 40968, 41067, 
    41166, 41264, 41363, 41462, 41561, 41659, 41758, 41857, 41956, 42054, 
    42153, 42252, 42350, 42449, 42548, 42646, 42745, 42844, 42942, 43041, 
    43140, 43238, 43337, 43436, 43534, 43633, 43732, 43830, 43929, 44028, 
    44126, 44225, 44324, 44422, 44521, 44619, 44718, 44817, 44915, 45014, 
    45112, 45211, 45310, 45408, 45507, 45605, 45704, 45802, 45901, 46000, 
    46098, 46197, 46295, 46394, 46492, 46591, 46689, 46788, 46886, 46985, 
    47084, 47182, 47281, 47379, 47478, 47576, 47675, 47773, 47872, 47970, 
    48069, 48167, 48266, 48364, 48462, 48561, 48659, 48758, 48856, 48955, 
    49053, 49152, 49250, 49349, 49447, 49545, 49644, 49742, 49841, 49939, 
    50038, 50136, 50234, 50333, 50431, 50530, 50628, 50726, 50825, 50923, 
    51022, 51120, 51218, 51317, 51415, 51513, 51612, 51710, 51809, 51907, 
    52005, 52104, 52202, 52300, 52399, 52497, 52595, 52694, 52792, 52890, 
    52989, 53087, 53185, 53283, 53382, 53480, 53578, 53677, 53775, 53873, 
    53972, 54070, 54168, 54266, 54365, 54463, 54561, 54659, 54758, 54856, 
    54954, 55052, 55151, 55249, 55347, 55445, 55544, 55642, 55740, 55838, 
    55937, 56035, 56133, 56231, 56329, 56428, 56526, 56624, 56722, 56820, 
    56919, 57017, 57115, 57213, 57311, 57409, 57508, 57606, 57704, 57802, 
    57900, 57998, 58097, 58195, 58293, 58391, 58489, 58587, 58685, 58784, 
    58882, 58980, 59078, 59176, 59274, 59372, 59470, 59568, 59666, 59765, 
    59863, 59961, 60059, 60157, 60255, 60353, 60451, 60549, 60647, 60745, 
    60843, 60941, 61040, 61138, 61236, 61334, 61432, 61530, 61628, 61726, 
    61824, 61922, 62020, 62118, 62216, 62314, 62412, 62510, 62608, 62706, 
    62804, 62902, 63000, 63098, 63196, 63294, 63392, 63490, 63588, 63686, 
    63784, 63882, 63980, 64077, 64175, 64273, 64371, 64469, 64567, 64665, 
    64763, 64861, 64959, 65057, 65155, 65253, 65351, 65448, 65546, 65644, 
    65742, 65840, 65938, 66036, 66134, 66232, 66330, 66427, 66525, 66623, 
    66721, 66819, 66917, 67015, 67112, 67210, 67308, 67406, 67504, 67602, 
    67700, 67797, 67895, 67993, 68091, 68189, 68286, 68384, 68482, 68580, 
    68678, 68775, 68873, 68971, 69069, 69167, 69264, 69362, 69460, 69558, 
    69656, 69753, 69851, 69949, 70047, 70144, 70242, 70340, 70438, 70535, 
    70633, 70731, 70829, 70926, 71024, 71122, 71219, 71317, 71415, 71513, 
    71610, 71708, 71806, 71903, 72001, 72099, 72197, 72294, 72392, 72490, 
    72587, 72685, 72783, 72880, 72978, 73076, 73173, 73271, 73369, 73466, 
    73564, 73662, 73759, 73857, 73954, 74052, 74150, 74247, 74345, 74442, 
    74540, 74638, 74735, 74833, 74931, 75028, 75126, 75223, 75321, 75419, 
    75516, 75614, 75711, 75809, 75906, 76004, 76102, 76199, 76297, 76394, 
    76492, 76589, 76687, 76784, 76882, 76979, 77077, 77175, 77272, 77370, 
    77467, 77565, 77662, 77760, 77857, 77955, 78052, 78150, 78247, 78345, 
    78442, 78540, 78637, 78735, 78832, 78930, 79027, 79124, 79222, 79319, 
    79417, 79514, 79612, 79709, 79807, 79904, 80001, 80099, 80196, 80294, 
    80391, 80489, 80586, 80683, 80781, 80878, 80976, 81073, 81170, 81268, 
    81365, 81463, 81560, 81657, 81755, 81852, 81950, 82047, 82144, 82242, 
    82339, 82436, 82534, 82631, 82728, 82826, 82923, 83020, 83118, 83215, 
    83312, 83410, 83507, 83604, 83702, 83799, 83896, 83994, 84091, 84188, 
    84286, 84383, 84480, 84577, 84675, 84772, 84869, 84967, 85064, 85161, 
    85258, 85356, 85453, 85550, 85647, 85745, 85842, 85939, 86036, 86134, 
    86231, 86328, 86425, 86523, 86620, 86717, 86814, 86911, 87009, 87106, 
    87203, 87300, 87398, 87495, 87592, 87689, 87786, 87883, 87981, 88078, 
    88175, 88272, 88369, 88466, 88564, 88661, 88758, 88855, 88952, 89049, 
    89147, 89244, 89341, 89438, 89535, 89632, 89729, 89826, 89924, 90021, 
    90118, 90215, 90312, 90409, 90506, 90603, 90700, 90797, 90895, 90992, 
    91089, 91186, 91283, 91380, 91477, 91574, 91671, 91768, 91865, 91962, 
    92059, 92156, 92253, 92351, 92448, 92545, 92642, 92739, 92836, 92933, 
    93030, 93127, 93224, 93321, 93418, 93515, 93612, 93709, 93806, 93903, 
    94000, 94097, 94194, 94291, 94388, 94485, 94581, 94678, 94775, 94872, 
    94969, 95066, 95163, 95260, 95357, 95454, 95551, 95648, 95745, 95842, 
    95939, 96036, 96132, 96229, 96326, 96423, 96520, 96617, 96714, 96811, 
    96908, 97005, 97102, 97198, 97295, 97392, 97489, 97586, 97683, 97780, 
    97876, 97973, 98070, 98167, 98264, 98361, 98458 ;

 refrac =
  27.079, 26.642, 26.213, 25.788, 25.366, 24.945, 24.527, 24.11, 23.695, 
    23.283, 22.879, 22.49, 22.119, 21.768, 21.432, 21.11, 20.797, 20.49, 
    20.186, 19.886, 19.588, 19.292, 18.998, 18.707, 18.419, 18.134, 17.852, 
    17.575, 17.302, 17.032, 16.765, 16.501, 16.253, 16.007, 15.762, 15.518, 
    15.273, 15.029, 14.786, 14.544, 14.305, 14.071, 13.842, 13.62, 13.405, 
    13.196, 12.995, 12.799, 12.608, 12.42, 12.235, 12.051, 11.867, 11.681, 
    11.495, 11.306, 11.117, 10.927, 10.738, 10.55, 10.364, 10.182, 10.005, 
    9.8329, 9.6664, 9.5058, 9.351, 9.2017, 9.0572, 8.9171, 8.7806, 8.6472, 
    8.5164, 8.3881, 8.262, 8.138, 8.0162, 7.8964, 7.7787, 7.6631, 7.5494, 
    7.4376, 7.3276, 7.2194, 7.1127, 7.0075, 6.9037, 6.801, 6.6995, 6.5991, 
    6.4999, 6.402, 6.3053, 6.2099, 6.1157, 6.0225, 5.9304, 5.8392, 5.749, 
    5.6597, 5.5716, 5.4847, 5.3992, 5.3152, 5.2328, 5.1521, 5.0732, 4.9962, 
    4.921, 4.8477, 4.7759, 4.7056, 4.6364, 4.5681, 4.5006, 4.4339, 4.3679, 
    4.3028, 4.2385, 4.1752, 4.1127, 4.0512, 3.9907, 3.9311, 3.8724, 3.8146, 
    3.7575, 3.701, 3.6449, 3.5892, 3.5339, 3.4791, 3.4249, 3.3716, 3.3191, 
    3.2676, 3.217, 3.1673, 3.1183, 3.0701, 3.0228, 2.9765, 2.9313, 2.8873, 
    2.8446, 2.8032, 2.7628, 2.7234, 2.6847, 2.6467, 2.6091, 2.5719, 2.535, 
    2.4983, 2.4618, 2.4256, 2.3898, 2.3546, 2.3199, 2.2859, 2.2527, 2.2201, 
    2.1881, 2.1567, 2.1257, 2.0951, 2.0649, 2.0351, 2.0056, 1.9766, 1.9478, 
    1.9194, 1.8914, 1.8636, 1.8361, 1.8089, 1.782, 1.7555, 1.7294, 1.7036, 
    1.6783, 1.6533, 1.6286, 1.6042, 1.58, 1.5561, 1.5325, 1.5093, 1.4864, 
    1.4639, 1.4418, 1.42, 1.3984, 1.3771, 1.356, 1.3353, 1.3148, 1.2947, 
    1.2749, 1.2556, 1.2366, 1.2179, 1.1997, 1.1819, 1.1644, 1.1471, 1.1302, 
    1.1135, 1.0969, 1.0806, 1.0644, 1.0484, 1.0328, 1.0174, 1.0025, 0.98808, 
    0.97415, 0.96071, 0.94772, 0.93512, 0.92283, 0.91079, 0.89891, 0.88711, 
    0.87532, 0.86352, 0.85167, 0.83981, 0.82796, 0.81617, 0.8045, 0.79302, 
    0.78177, 0.7708, 0.76009, 0.74961, 0.73935, 0.72929, 0.71942, 0.70973, 
    0.70021, 0.69086, 0.68169, 0.67269, 0.66387, 0.65525, 0.64681, 0.63852, 
    0.63034, 0.62223, 0.61415, 0.60608, 0.59801, 0.58994, 0.58187, 0.57387, 
    0.56599, 0.55828, 0.5508, 0.54356, 0.53655, 0.52974, 0.52309, 0.51656, 
    0.51011, 0.50371, 0.49732, 0.49092, 0.4845, 0.47807, 0.47164, 0.46528, 
    0.45902, 0.45295, 0.44714, 0.4416, 0.43632, 0.43122, 0.42618, 0.42108, 
    0.41585, 0.41044, 0.40489, 0.39925, 0.39364, 0.38817, 0.38298, 0.37815, 
    0.37375, 0.36977, 0.36613, 0.36271, 0.35933, 0.35581, 0.35198, 0.34772, 
    0.343, 0.33787, 0.33245, 0.32692, 0.32149, 0.31636, 0.31167, 0.30749, 
    0.30382, 0.30055, 0.29755, 0.29468, 0.2918, 0.28887, 0.28586, 0.28281, 
    0.27975, 0.27673, 0.27377, 0.27086, 0.26797, 0.26508, 0.26215, 0.25915, 
    0.25605, 0.25285, 0.24958, 0.24626, 0.24293, 0.23962, 0.23637, 0.23319, 
    0.23008, 0.22703, 0.22402, 0.22103, 0.21804, 0.21506, 0.21213, 0.20928, 
    0.20656, 0.204, 0.20162, 0.19941, 0.19732, 0.1953, 0.19328, 0.19119, 
    0.18902, 0.18676, 0.18445, 0.18211, 0.17979, 0.17752, 0.17533, 0.17321, 
    0.17115, 0.16913, 0.16713, 0.16512, 0.16308, 0.161, 0.15889, 0.15677, 
    0.15467, 0.15262, 0.15063, 0.14873, 0.1469, 0.14515, 0.14345, 0.14179, 
    0.14013, 0.13846, 0.13676, 0.13504, 0.13334, 0.13167, 0.13006, 0.12851, 
    0.12703, 0.12561, 0.12422, 0.12285, 0.1215, 0.12017, 0.11886, 0.11758, 
    0.11632, 0.11508, 0.11384, 0.11259, 0.11132, 0.11001, 0.10868, 0.10732, 
    0.10595, 0.10456, 0.10318, 0.10181, 0.10048, 0.099173, 0.097911, 
    0.096685, 0.095488, 0.094312, 0.09315, 0.091998, 0.090853, 0.08971, 
    0.088567, 0.087423, 0.086279, 0.085138, 0.084003, 0.082877, 0.081763, 
    0.080665, 0.079589, 0.078545, 0.07754, 0.07658, 0.075667, 0.074797, 
    0.073962, 0.073148, 0.072341, 0.071528, 0.0707, 0.069855, 0.068999, 
    0.068138, 0.067282, 0.066436, 0.065602, 0.064777, 0.063957, 0.063136, 
    0.062309, 0.061473, 0.060628, 0.059777, 0.058925, 0.058084, 0.057266, 
    0.056479, 0.055734, 0.055036, 0.054385, 0.053774, 0.05319, 0.052617, 
    0.052037, 0.051438, 0.050812, 0.050161, 0.049491, 0.04881, 0.048131, 
    0.047466, 0.046823, 0.046209, 0.045625, 0.045066, 0.044523, 0.043984, 
    0.043439, 0.042879, 0.042301, 0.041708, 0.041106, 0.040504, 0.039909, 
    0.03933, 0.038774, 0.038244, 0.037737, 0.037251, 0.03678, 0.036316, 
    0.035853, 0.035388, 0.034918, 0.034445, 0.033974, 0.033508, 0.03305, 
    0.032602, 0.032166, 0.031738, 0.031319, 0.030905, 0.030495, 0.030085, 
    0.029674, 0.029259, 0.028842, 0.028425, 0.028012, 0.027607, 0.027213, 
    0.026831, 0.02646, 0.026099, 0.025745, 0.025396, 0.02505, 0.024707, 
    0.024367, 0.024031, 0.0237, 0.023373, 0.023049, 0.022728, 0.02241, 
    0.022094, 0.021781, 0.021471, 0.021163, 0.020859, 0.020558, 0.020262, 
    0.019971, 0.019687, 0.019409, 0.019137, 0.01887, 0.018608, 0.018349, 
    0.018092, 0.017836, 0.017582, 0.01733, 0.017081, 0.016836, 0.016596, 
    0.016362, 0.016133, 0.015907, 0.015685, 0.015464, 0.015244, 0.015026, 
    0.014809, 0.014594, 0.014381, 0.014171, 0.013965, 0.013762, 0.013562, 
    0.013366, 0.013172, 0.01298, 0.01279, 0.012603, 0.012418, 0.012235, 
    0.012054, 0.011875, 0.0117, 0.011528, 0.011359, 0.011192, 0.011028, 
    0.010867, 0.010707, 0.01055, 0.010394, 0.01024, 0.010088, 0.0099378, 
    0.0097901, 0.0096446, 0.0095011, 0.0093595, 0.0092194, 0.009081, 
    0.0089448, 0.0088103, 0.0086776, 0.0085467, 0.0084176, 0.0082901, 
    0.0081644, 0.0080403, 0.0079179, 0.0077971, 0.0076779, 0.0075603, 
    0.0074443, 0.0073298, 0.0072169, 0.0071055, 0.0069955, 0.0068871, 
    0.0067801, 0.0066745, 0.0065703, 0.0064676, 0.0063662, 0.0062662, 
    0.0061676, 0.0060703, 0.0059743, 0.0058796, 0.0057862, 0.005694, 
    0.0056031, 0.0055135, 0.0054251, 0.0053379, 0.0052518, 0.005167, 
    0.0050833, 0.0050008, 0.0049194, 0.0048392, 0.0047601, 0.004682, 
    0.0046051, 0.0045292, 0.0044544, 0.0043806, 0.0043079, 0.0042362, 
    0.0041655, 0.0040958, 0.0040271, 0.0039594, 0.0038926, 0.0038268, 
    0.003762, 0.0036981, 0.0036351, 0.003573, 0.0035118, 0.0034515, 
    0.0033921, 0.0033335, 0.0032759, 0.003219, 0.0031631, 0.0031079, 
    0.0030536, 0.003, 0.0029473, 0.0028954, 0.0028442, 0.0027939, 0.0027443, 
    0.0026954, 0.0026473, 0.0025999, 0.0025533, 0.0025074, 0.0024622, 
    0.0024177, 0.0023739, 0.0023308, 0.0022884, 0.0022466, 0.0022055, 
    0.0021651, 0.0021253, 0.0020861, 0.0020476, 0.0020097, 0.0019724, 
    0.0019357, 0.0018996, 0.0018641, 0.0018292, 0.0017948, 0.0017611, 
    0.0017279, 0.0016952, 0.0016631, 0.0016316, 0.0016005, 0.00157, 
    0.0015401, 0.0015106, 0.0014816, 0.0014531, 0.0014252, 0.0013977, 
    0.0013707, 0.0013441, 0.0013181, 0.0012924, 0.0012673, 0.0012426, 
    0.0012183, 0.0011944, 0.001171, 0.001148, 0.0011254, 0.0011032, 
    0.0010815, 0.0010601, 0.0010391, 0.0010185, 0.00099827, 0.00097842, 
    0.00095894, 0.00093981, 0.00092104, 0.00090263, 0.00088455, 0.00086682, 
    0.00084942, 0.00083235, 0.00081561, 0.00079918, 0.00078307, 0.00076726, 
    0.00075176, 0.00073655, 0.00072164, 0.00070702, 0.00069268, 0.00067862, 
    0.00066483, 0.00065131, 0.00063806, 0.00062507, 0.00061233, 0.00059985, 
    0.00058761, 0.00057561, 0.00056386, 0.00055233, 0.00054104, 0.00052997, 
    0.00051913, 0.0005085, 0.00049809, 0.00048789, 0.00047789, 0.0004681, 
    0.00045851, 0.00044911, 0.0004399, 0.00043088, 0.00042204, 0.00041339, 
    0.00040491, 0.00039661, 0.00038848, 0.00038051, 0.00037271, 0.00036508, 
    0.0003576, 0.00035027, 0.0003431, 0.00033608, 0.0003292, 0.00032246, 
    0.00031587, 0.00030942, 0.0003031, 0.00029691, 0.00029085, 0.00028492, 
    0.00027911, 0.00027343, 0.00026786, 0.00026242, 0.00025708, 0.00025186, 
    0.00024675, 0.00024175, 0.00023685, 0.00023206, 0.00022737, 0.00022278, 
    0.00021828, 0.00021388, 0.00020958, 0.00020536, 0.00020124, 0.0001972, 
    0.00019325, 0.00018938, 0.00018559, 0.00018189, 0.00017826, 0.00017471, 
    0.00017124, 0.00016783, 0.00016451, 0.00016125, 0.00015806, 0.00015494, 
    0.00015188, 0.00014889, 0.00014597, 0.0001431, 0.0001403, 0.00013755, 
    0.00013487, 0.00013224, 0.00012966, 0.00012714, 0.00012468, 0.00012226, 
    0.0001199, 0.00011759, 0.00011532, 0.00011311, 0.00011094, 0.00010881, 
    0.00010673, 0.00010469, 0.0001027, 0.00010075, 9.8838e-05, 9.6967e-05, 
    9.5135e-05, 9.3341e-05, 9.1585e-05,
  27.079, 26.642, 26.213, 25.788, 25.366, 24.945, 24.527, 24.11, 23.695, 
    23.283, 22.879, 22.49, 22.119, 21.768, 21.432, 21.11, 20.797, 20.49, 
    20.186, 19.886, 19.588, 19.292, 18.998, 18.707, 18.419, 18.134, 17.852, 
    17.575, 17.302, 17.032, 16.765, 16.501, 16.253, 16.007, 15.762, 15.518, 
    15.273, 15.029, 14.786, 14.544, 14.305, 14.071, 13.842, 13.62, 13.405, 
    13.196, 12.995, 12.799, 12.608, 12.42, 12.235, 12.051, 11.867, 11.681, 
    11.495, 11.306, 11.117, 10.927, 10.738, 10.55, 10.364, 10.182, 10.005, 
    9.8329, 9.6664, 9.5058, 9.351, 9.2017, 9.0572, 8.9171, 8.7806, 8.6472, 
    8.5164, 8.3881, 8.262, 8.138, 8.0162, 7.8964, 7.7787, 7.6631, 7.5494, 
    7.4376, 7.3276, 7.2194, 7.1127, 7.0075, 6.9037, 6.801, 6.6995, 6.5991, 
    6.4999, 6.402, 6.3053, 6.2099, 6.1157, 6.0225, 5.9304, 5.8392, 5.749, 
    5.6597, 5.5716, 5.4847, 5.3992, 5.3152, 5.2328, 5.1521, 5.0732, 4.9962, 
    4.921, 4.8477, 4.7759, 4.7056, 4.6364, 4.5681, 4.5006, 4.4339, 4.3679, 
    4.3028, 4.2385, 4.1752, 4.1127, 4.0512, 3.9907, 3.9311, 3.8724, 3.8146, 
    3.7575, 3.701, 3.6449, 3.5892, 3.5339, 3.4791, 3.4249, 3.3716, 3.3191, 
    3.2676, 3.217, 3.1673, 3.1183, 3.0701, 3.0228, 2.9765, 2.9313, 2.8873, 
    2.8446, 2.8032, 2.7628, 2.7234, 2.6847, 2.6467, 2.6091, 2.5719, 2.535, 
    2.4983, 2.4618, 2.4256, 2.3898, 2.3546, 2.3199, 2.2859, 2.2527, 2.2201, 
    2.1881, 2.1567, 2.1257, 2.0951, 2.0649, 2.0351, 2.0056, 1.9766, 1.9478, 
    1.9194, 1.8914, 1.8636, 1.8361, 1.8089, 1.782, 1.7555, 1.7294, 1.7036, 
    1.6783, 1.6533, 1.6286, 1.6042, 1.58, 1.5561, 1.5325, 1.5093, 1.4864, 
    1.4639, 1.4418, 1.42, 1.3984, 1.3771, 1.356, 1.3353, 1.3148, 1.2947, 
    1.2749, 1.2556, 1.2366, 1.2179, 1.1997, 1.1819, 1.1644, 1.1471, 1.1302, 
    1.1135, 1.0969, 1.0806, 1.0644, 1.0484, 1.0328, 1.0174, 1.0025, 0.98808, 
    0.97415, 0.96071, 0.94772, 0.93512, 0.92283, 0.91079, 0.89891, 0.88711, 
    0.87532, 0.86352, 0.85167, 0.83981, 0.82796, 0.81617, 0.8045, 0.79302, 
    0.78177, 0.7708, 0.76009, 0.74961, 0.73935, 0.72929, 0.71942, 0.70973, 
    0.70021, 0.69086, 0.68169, 0.67269, 0.66387, 0.65525, 0.64681, 0.63852, 
    0.63034, 0.62223, 0.61415, 0.60608, 0.59801, 0.58994, 0.58187, 0.57387, 
    0.56599, 0.55828, 0.5508, 0.54356, 0.53655, 0.52974, 0.52309, 0.51656, 
    0.51011, 0.50371, 0.49732, 0.49092, 0.4845, 0.47807, 0.47164, 0.46528, 
    0.45902, 0.45295, 0.44714, 0.4416, 0.43632, 0.43122, 0.42618, 0.42108, 
    0.41585, 0.41044, 0.40489, 0.39925, 0.39364, 0.38817, 0.38298, 0.37815, 
    0.37375, 0.36977, 0.36613, 0.36271, 0.35933, 0.35581, 0.35198, 0.34772, 
    0.343, 0.33787, 0.33245, 0.32692, 0.32149, 0.31636, 0.31167, 0.30749, 
    0.30382, 0.30055, 0.29755, 0.29468, 0.2918, 0.28887, 0.28586, 0.28281, 
    0.27975, 0.27673, 0.27377, 0.27086, 0.26797, 0.26508, 0.26215, 0.25915, 
    0.25605, 0.25285, 0.24958, 0.24626, 0.24293, 0.23962, 0.23637, 0.23319, 
    0.23008, 0.22703, 0.22402, 0.22103, 0.21804, 0.21506, 0.21213, 0.20928, 
    0.20656, 0.204, 0.20162, 0.19941, 0.19732, 0.1953, 0.19328, 0.19119, 
    0.18902, 0.18676, 0.18445, 0.18211, 0.17979, 0.17752, 0.17533, 0.17321, 
    0.17115, 0.16913, 0.16713, 0.16512, 0.16308, 0.161, 0.15889, 0.15677, 
    0.15467, 0.15262, 0.15063, 0.14873, 0.1469, 0.14515, 0.14345, 0.14179, 
    0.14013, 0.13846, 0.13676, 0.13504, 0.13334, 0.13167, 0.13006, 0.12851, 
    0.12703, 0.12561, 0.12422, 0.12285, 0.1215, 0.12017, 0.11886, 0.11758, 
    0.11632, 0.11508, 0.11384, 0.11259, 0.11132, 0.11001, 0.10868, 0.10732, 
    0.10595, 0.10456, 0.10318, 0.10181, 0.10048, 0.099173, 0.097911, 
    0.096685, 0.095488, 0.094312, 0.09315, 0.091998, 0.090853, 0.08971, 
    0.088567, 0.087423, 0.086279, 0.085138, 0.084003, 0.082877, 0.081763, 
    0.080665, 0.079589, 0.078545, 0.07754, 0.07658, 0.075667, 0.074797, 
    0.073962, 0.073148, 0.072341, 0.071528, 0.0707, 0.069855, 0.068999, 
    0.068138, 0.067282, 0.066436, 0.065602, 0.064777, 0.063957, 0.063136, 
    0.062309, 0.061473, 0.060628, 0.059777, 0.058925, 0.058084, 0.057266, 
    0.056479, 0.055734, 0.055036, 0.054385, 0.053774, 0.05319, 0.052617, 
    0.052037, 0.051438, 0.050812, 0.050161, 0.049491, 0.04881, 0.048131, 
    0.047466, 0.046823, 0.046209, 0.045625, 0.045066, 0.044523, 0.043984, 
    0.043439, 0.042879, 0.042301, 0.041708, 0.041106, 0.040504, 0.039909, 
    0.03933, 0.038774, 0.038244, 0.037737, 0.037251, 0.03678, 0.036316, 
    0.035853, 0.035388, 0.034918, 0.034445, 0.033974, 0.033508, 0.03305, 
    0.032602, 0.032166, 0.031738, 0.031319, 0.030905, 0.030495, 0.030085, 
    0.029674, 0.029259, 0.028842, 0.028425, 0.028012, 0.027607, 0.027213, 
    0.026831, 0.02646, 0.026099, 0.025745, 0.025396, 0.02505, 0.024707, 
    0.024367, 0.024031, 0.0237, 0.023373, 0.023049, 0.022728, 0.02241, 
    0.022094, 0.021781, 0.021471, 0.021163, 0.020859, 0.020558, 0.020262, 
    0.019971, 0.019687, 0.019409, 0.019137, 0.01887, 0.018608, 0.018349, 
    0.018092, 0.017836, 0.017582, 0.01733, 0.017081, 0.016836, 0.016596, 
    0.016362, 0.016133, 0.015907, 0.015685, 0.015464, 0.015244, 0.015026, 
    0.014809, 0.014594, 0.014381, 0.014171, 0.013965, 0.013762, 0.013562, 
    0.013366, 0.013172, 0.01298, 0.01279, 0.012603, 0.012418, 0.012235, 
    0.012054, 0.011875, 0.0117, 0.011528, 0.011359, 0.011192, 0.011028, 
    0.010867, 0.010707, 0.01055, 0.010394, 0.01024, 0.010088, 0.0099378, 
    0.0097901, 0.0096446, 0.0095011, 0.0093595, 0.0092194, 0.009081, 
    0.0089448, 0.0088103, 0.0086776, 0.0085467, 0.0084176, 0.0082901, 
    0.0081644, 0.0080403, 0.0079179, 0.0077971, 0.0076779, 0.0075603, 
    0.0074443, 0.0073298, 0.0072169, 0.0071055, 0.0069955, 0.0068871, 
    0.0067801, 0.0066745, 0.0065703, 0.0064676, 0.0063662, 0.0062662, 
    0.0061676, 0.0060703, 0.0059743, 0.0058796, 0.0057862, 0.005694, 
    0.0056031, 0.0055135, 0.0054251, 0.0053379, 0.0052518, 0.005167, 
    0.0050833, 0.0050008, 0.0049194, 0.0048392, 0.0047601, 0.004682, 
    0.0046051, 0.0045292, 0.0044544, 0.0043806, 0.0043079, 0.0042362, 
    0.0041655, 0.0040958, 0.0040271, 0.0039594, 0.0038926, 0.0038268, 
    0.003762, 0.0036981, 0.0036351, 0.003573, 0.0035118, 0.0034515, 
    0.0033921, 0.0033335, 0.0032759, 0.003219, 0.0031631, 0.0031079, 
    0.0030536, 0.003, 0.0029473, 0.0028954, 0.0028442, 0.0027939, 0.0027443, 
    0.0026954, 0.0026473, 0.0025999, 0.0025533, 0.0025074, 0.0024622, 
    0.0024177, 0.0023739, 0.0023308, 0.0022884, 0.0022466, 0.0022055, 
    0.0021651, 0.0021253, 0.0020861, 0.0020476, 0.0020097, 0.0019724, 
    0.0019357, 0.0018996, 0.0018641, 0.0018292, 0.0017948, 0.0017611, 
    0.0017279, 0.0016952, 0.0016631, 0.0016316, 0.0016005, 0.00157, 
    0.0015401, 0.0015106, 0.0014816, 0.0014531, 0.0014252, 0.0013977, 
    0.0013707, 0.0013441, 0.0013181, 0.0012924, 0.0012673, 0.0012426, 
    0.0012183, 0.0011944, 0.001171, 0.001148, 0.0011254, 0.0011032, 
    0.0010815, 0.0010601, 0.0010391, 0.0010185, 0.00099827, 0.00097842, 
    0.00095894, 0.00093981, 0.00092104, 0.00090263, 0.00088455, 0.00086682, 
    0.00084942, 0.00083235, 0.00081561, 0.00079918, 0.00078307, 0.00076726, 
    0.00075176, 0.00073655, 0.00072164, 0.00070702, 0.00069268, 0.00067862, 
    0.00066483, 0.00065131, 0.00063806, 0.00062507, 0.00061233, 0.00059985, 
    0.00058761, 0.00057561, 0.00056386, 0.00055233, 0.00054104, 0.00052997, 
    0.00051913, 0.0005085, 0.00049809, 0.00048789, 0.00047789, 0.0004681, 
    0.00045851, 0.00044911, 0.0004399, 0.00043088, 0.00042204, 0.00041339, 
    0.00040491, 0.00039661, 0.00038848, 0.00038051, 0.00037271, 0.00036508, 
    0.0003576, 0.00035027, 0.0003431, 0.00033608, 0.0003292, 0.00032246, 
    0.00031587, 0.00030942, 0.0003031, 0.00029691, 0.00029085, 0.00028492, 
    0.00027911, 0.00027343, 0.00026786, 0.00026242, 0.00025708, 0.00025186, 
    0.00024675, 0.00024175, 0.00023685, 0.00023206, 0.00022737, 0.00022278, 
    0.00021828, 0.00021388, 0.00020958, 0.00020536, 0.00020124, 0.0001972, 
    0.00019325, 0.00018938, 0.00018559, 0.00018189, 0.00017826, 0.00017471, 
    0.00017124, 0.00016783, 0.00016451, 0.00016125, 0.00015806, 0.00015494, 
    0.00015188, 0.00014889, 0.00014597, 0.0001431, 0.0001403, 0.00013755, 
    0.00013487, 0.00013224, 0.00012966, 0.00012714, 0.00012468, 0.00012226, 
    0.0001199, 0.00011759, 0.00011532, 0.00011311, 0.00011094, 0.00010881, 
    0.00010673, 0.00010469, 0.0001027, 0.00010075, 9.8838e-05, 9.6967e-05, 
    9.5135e-05, 9.3341e-05, 9.1585e-05 ;

 refrac_sigma =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 refrac_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07 ;

 dry_temp =
  250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250,
  250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250 ;

 dry_temp_sigma =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07 ;

 dry_temp_qual =
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07,
  -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, -9.9999e+07, 
    -9.9999e+07, -9.9999e+07 ;
}
